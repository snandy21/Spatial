`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif

module RetimeWrapper(
  input   clock,
  input   reset,
  input   io_flow,
  input   io_in,
  output  io_out
);
  wire  sr_out;
  wire  sr_in;
  wire  sr_flow;
  wire  sr_reset;
  wire  sr_clock;
  RetimeShiftRegister #(.WIDTH(1), .STAGES(1)) sr (
    .out(sr_out),
    .in(sr_in),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out;
  assign sr_in = io_in;
  assign sr_flow = io_flow;
  assign sr_reset = reset;
  assign sr_clock = clock;
endmodule
module FF(
  input        clock,
  input        reset,
  input  [7:0] io_input_0_data,
  input        io_input_0_enable,
  input        io_input_0_reset,
  output [7:0] io_output_data
);
  reg [7:0] ff;
  reg [31:0] _RAND_0;
  wire [7:0] _T_7;
  wire [7:0] _T_8;
  wire [7:0] _T_9;
  assign _T_7 = io_input_0_enable ? io_input_0_data : ff;
  assign _T_8 = io_input_0_reset ? 8'h0 : _T_7;
  assign _T_9 = io_input_0_reset ? 8'h0 : ff;
  assign io_output_data = _T_9;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  ff = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 8'h0;
    end else begin
      if (io_input_0_reset) begin
        ff <= 8'h0;
      end else begin
        if (io_input_0_enable) begin
          ff <= io_input_0_data;
        end
      end
    end
  end
endmodule
module SingleCounter(
  input        clock,
  input        reset,
  input  [7:0] io_input_stop,
  input        io_input_reset,
  input        io_input_enable,
  output       io_output_done
);
  wire  FF_clock;
  wire  FF_reset;
  wire [7:0] FF_io_input_0_data;
  wire  FF_io_input_0_enable;
  wire  FF_io_input_0_reset;
  wire [7:0] FF_io_output_data;
  wire [7:0] _T_21;
  wire [8:0] _T_23;
  wire [7:0] _T_24;
  wire [7:0] _T_25;
  wire  _T_28;
  wire [7:0] _T_38;
  wire [7:0] _T_41;
  wire [7:0] _T_42;
  wire [7:0] _T_43;
  wire  _T_47;
  FF FF (
    .clock(FF_clock),
    .reset(FF_reset),
    .io_input_0_data(FF_io_input_0_data),
    .io_input_0_enable(FF_io_input_0_enable),
    .io_input_0_reset(FF_io_input_0_reset),
    .io_output_data(FF_io_output_data)
  );
  assign _T_21 = $signed(FF_io_output_data);
  assign _T_23 = $signed(_T_21) + $signed(8'sh1);
  assign _T_24 = _T_23[7:0];
  assign _T_25 = $signed(_T_24);
  assign _T_28 = $signed(_T_25) >= $signed(io_input_stop);
  assign _T_38 = $unsigned(_T_21);
  assign _T_41 = $unsigned(_T_25);
  assign _T_42 = _T_28 ? _T_38 : _T_41;
  assign _T_43 = io_input_reset ? 8'h0 : _T_42;
  assign _T_47 = io_input_enable & _T_28;
  assign io_output_done = _T_47;
  assign FF_io_input_0_data = _T_43;
  assign FF_io_input_0_enable = io_input_enable;
  assign FF_io_input_0_reset = io_input_reset;
  assign FF_clock = clock;
  assign FF_reset = reset;
endmodule
module SRFF(
  input   clock,
  input   reset,
  input   io_input_set,
  input   io_input_reset,
  input   io_input_asyn_reset,
  output  io_output_data
);
  reg  _T_8;
  reg [31:0] _RAND_0;
  wire  _T_12;
  wire  _T_13;
  wire  _T_14;
  wire  _T_16;
  assign _T_12 = io_input_reset ? 1'h0 : _T_8;
  assign _T_13 = io_input_set ? 1'h1 : _T_12;
  assign _T_14 = io_input_asyn_reset ? 1'h0 : _T_13;
  assign _T_16 = io_input_asyn_reset ? 1'h0 : _T_8;
  assign io_output_data = _T_16;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_8 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_8 <= 1'h0;
    end else begin
      if (io_input_asyn_reset) begin
        _T_8 <= 1'h0;
      end else begin
        if (io_input_set) begin
          _T_8 <= 1'h1;
        end else begin
          if (io_input_reset) begin
            _T_8 <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module FF_1(
  input         clock,
  input         reset,
  input  [31:0] io_input_0_data,
  input  [31:0] io_input_0_init,
  input         io_input_0_enable,
  input         io_input_0_reset,
  output [31:0] io_output_data
);
  reg [31:0] ff;
  reg [31:0] _RAND_0;
  wire [31:0] _T_7;
  wire [31:0] _T_8;
  wire [31:0] _T_9;
  assign _T_7 = io_input_0_enable ? io_input_0_data : ff;
  assign _T_8 = io_input_0_reset ? io_input_0_init : _T_7;
  assign _T_9 = io_input_0_reset ? io_input_0_init : ff;
  assign io_output_data = _T_9;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  ff = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= io_input_0_init;
    end else begin
      if (io_input_0_reset) begin
        ff <= io_input_0_init;
      end else begin
        if (io_input_0_enable) begin
          ff <= io_input_0_data;
        end
      end
    end
  end
endmodule
module RetimeWrapper_6(
  input         clock,
  input         reset,
  input  [31:0] io_in,
  output [31:0] io_out
);
  wire [31:0] sr_out;
  wire [31:0] sr_in;
  wire  sr_flow;
  wire  sr_reset;
  wire  sr_clock;
  RetimeShiftRegister #(.WIDTH(32), .STAGES(1)) sr (
    .out(sr_out),
    .in(sr_in),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out;
  assign sr_in = io_in;
  assign sr_flow = 1'h1;
  assign sr_reset = reset;
  assign sr_clock = clock;
endmodule
module SingleCounter_1(
  input         clock,
  input         reset,
  input  [31:0] io_input_stop,
  input  [31:0] io_input_stride,
  input         io_input_reset,
  input         io_input_enable,
  input         io_input_saturate,
  output [31:0] io_output_count_0,
  output        io_output_done
);
  wire  FF_clock;
  wire  FF_reset;
  wire [31:0] FF_io_input_0_data;
  wire [31:0] FF_io_input_0_init;
  wire  FF_io_input_0_enable;
  wire  FF_io_input_0_reset;
  wire [31:0] FF_io_output_data;
  wire [31:0] _T_21;
  wire [32:0] _T_23;
  wire [31:0] _T_24;
  wire [31:0] _T_25;
  wire  _T_27;
  wire  _T_28;
  wire  _T_29;
  wire  _T_30;
  wire [31:0] _T_38;
  wire [31:0] _T_40;
  wire [31:0] _T_41;
  wire [31:0] _T_42;
  wire [31:0] _T_43;
  wire  _T_47;
  FF_1 FF (
    .clock(FF_clock),
    .reset(FF_reset),
    .io_input_0_data(FF_io_input_0_data),
    .io_input_0_init(FF_io_input_0_init),
    .io_input_0_enable(FF_io_input_0_enable),
    .io_input_0_reset(FF_io_input_0_reset),
    .io_output_data(FF_io_output_data)
  );
  assign _T_21 = $signed(FF_io_output_data);
  assign _T_23 = $signed(_T_21) + $signed(32'sh1);
  assign _T_24 = _T_23[31:0];
  assign _T_25 = $signed(_T_24);
  assign _T_27 = $signed(io_input_stride) >= $signed(32'sh0);
  assign _T_28 = $signed(_T_25) >= $signed(io_input_stop);
  assign _T_29 = $signed(_T_25) <= $signed(io_input_stop);
  assign _T_30 = _T_27 ? _T_28 : _T_29;
  assign _T_38 = $unsigned(_T_21);
  assign _T_40 = io_input_saturate ? _T_38 : 32'h0;
  assign _T_41 = $unsigned(_T_25);
  assign _T_42 = _T_30 ? _T_40 : _T_41;
  assign _T_43 = io_input_reset ? 32'h0 : _T_42;
  assign _T_47 = io_input_enable & _T_30;
  assign io_output_count_0 = _T_21;
  assign io_output_done = _T_47;
  assign FF_io_input_0_data = _T_43;
  assign FF_io_input_0_init = 32'h0;
  assign FF_io_input_0_enable = io_input_enable;
  assign FF_io_input_0_reset = io_input_reset;
  assign FF_clock = clock;
  assign FF_reset = reset;
endmodule
module Seqpipe(
  input   clock,
  input   reset,
  input   io_input_enable,
  input   io_input_stageDone_0,
  input   io_input_stageDone_1,
  input   io_input_stageMask_0,
  input   io_input_stageMask_1,
  input   io_input_rst,
  output  io_output_done,
  output  io_output_stageEnable_0,
  output  io_output_stageEnable_1,
  output  io_output_rst_en
);
  wire  SingleCounter_clock;
  wire  SingleCounter_reset;
  wire [7:0] SingleCounter_io_input_stop;
  wire  SingleCounter_io_input_reset;
  wire  SingleCounter_io_input_enable;
  wire  SingleCounter_io_output_done;
  wire  SRFF_clock;
  wire  SRFF_reset;
  wire  SRFF_io_input_set;
  wire  SRFF_io_input_reset;
  wire  SRFF_io_input_asyn_reset;
  wire  SRFF_io_output_data;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire  RetimeWrapper_io_flow;
  wire  RetimeWrapper_io_in;
  wire  RetimeWrapper_io_out;
  wire  _T_26;
  wire  RetimeWrapper_1_clock;
  wire  RetimeWrapper_1_reset;
  wire  RetimeWrapper_1_io_flow;
  wire  RetimeWrapper_1_io_in;
  wire  RetimeWrapper_1_io_out;
  wire  _T_30;
  wire  FF_clock;
  wire  FF_reset;
  wire [31:0] FF_io_input_0_data;
  wire [31:0] FF_io_input_0_init;
  wire  FF_io_input_0_enable;
  wire  FF_io_input_0_reset;
  wire [31:0] FF_io_output_data;
  wire  RetimeWrapper_2_clock;
  wire  RetimeWrapper_2_reset;
  wire  RetimeWrapper_2_io_flow;
  wire  RetimeWrapper_2_io_in;
  wire  RetimeWrapper_2_io_out;
  wire  _T_36;
  wire [31:0] _T_37;
  wire  _T_39;
  wire  _T_40;
  wire  _T_42;
  wire  RetimeWrapper_3_clock;
  wire  RetimeWrapper_3_reset;
  wire  RetimeWrapper_3_io_flow;
  wire  RetimeWrapper_3_io_in;
  wire  RetimeWrapper_3_io_out;
  wire  _T_46;
  wire  _T_47;
  wire [7:0] _T_51;
  wire  FF_1_clock;
  wire  FF_1_reset;
  wire [31:0] FF_1_io_input_0_data;
  wire [31:0] FF_1_io_input_0_init;
  wire  FF_1_io_input_0_enable;
  wire  FF_1_io_input_0_reset;
  wire [31:0] FF_1_io_output_data;
  wire  RetimeWrapper_4_clock;
  wire  RetimeWrapper_4_reset;
  wire  RetimeWrapper_4_io_flow;
  wire  RetimeWrapper_4_io_in;
  wire  RetimeWrapper_4_io_out;
  wire  _T_58;
  wire  RetimeWrapper_5_clock;
  wire  RetimeWrapper_5_reset;
  wire [31:0] RetimeWrapper_5_io_in;
  wire [31:0] RetimeWrapper_5_io_out;
  wire [31:0] _T_63;
  wire  SingleCounter_1_clock;
  wire  SingleCounter_1_reset;
  wire [31:0] SingleCounter_1_io_input_stop;
  wire [31:0] SingleCounter_1_io_input_stride;
  wire  SingleCounter_1_io_input_reset;
  wire  SingleCounter_1_io_input_enable;
  wire  SingleCounter_1_io_input_saturate;
  wire [31:0] SingleCounter_1_io_output_count_0;
  wire  SingleCounter_1_io_output_done;
  wire  _T_64;
  wire [31:0] _T_66;
  wire  RetimeWrapper_6_clock;
  wire  RetimeWrapper_6_reset;
  wire  RetimeWrapper_6_io_flow;
  wire  RetimeWrapper_6_io_in;
  wire  RetimeWrapper_6_io_out;
  wire  _T_70;
  wire  _T_72;
  wire  _T_73;
  wire  RetimeWrapper_7_clock;
  wire  RetimeWrapper_7_reset;
  wire  RetimeWrapper_7_io_flow;
  wire  RetimeWrapper_7_io_in;
  wire  RetimeWrapper_7_io_out;
  wire  _T_79;
  wire [1:0] _T_91;
  wire [2:0] _T_92;
  wire  _T_96;
  wire  _T_98;
  wire  _T_99;
  wire  _T_101;
  wire  _T_102;
  wire [32:0] _T_104;
  wire [31:0] _T_105;
  wire [31:0] _T_106;
  wire [31:0] _T_107;
  wire  _T_109;
  wire  _T_110;
  wire  _T_111;
  wire  _T_112;
  wire [32:0] _T_114;
  wire [31:0] _T_115;
  wire [31:0] _T_116;
  wire [31:0] _T_117;
  wire [31:0] _T_118;
  wire [31:0] _GEN_0;
  wire  _T_120;
  wire [2:0] _GEN_1;
  wire [31:0] _GEN_2;
  wire [31:0] _GEN_3;
  wire [31:0] _GEN_4;
  wire [31:0] _GEN_5;
  wire [31:0] _GEN_6;
  wire [31:0] _GEN_8;
  wire  _T_144;
  SingleCounter SingleCounter (
    .clock(SingleCounter_clock),
    .reset(SingleCounter_reset),
    .io_input_stop(SingleCounter_io_input_stop),
    .io_input_reset(SingleCounter_io_input_reset),
    .io_input_enable(SingleCounter_io_input_enable),
    .io_output_done(SingleCounter_io_output_done)
  );
  SRFF SRFF (
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output_data(SRFF_io_output_data)
  );
  RetimeWrapper RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 (
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  FF_1 FF (
    .clock(FF_clock),
    .reset(FF_reset),
    .io_input_0_data(FF_io_input_0_data),
    .io_input_0_init(FF_io_input_0_init),
    .io_input_0_enable(FF_io_input_0_enable),
    .io_input_0_reset(FF_io_input_0_reset),
    .io_output_data(FF_io_output_data)
  );
  RetimeWrapper RetimeWrapper_2 (
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 (
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  FF_1 FF_1 (
    .clock(FF_1_clock),
    .reset(FF_1_reset),
    .io_input_0_data(FF_1_io_input_0_data),
    .io_input_0_init(FF_1_io_input_0_init),
    .io_input_0_enable(FF_1_io_input_0_enable),
    .io_input_0_reset(FF_1_io_input_0_reset),
    .io_output_data(FF_1_io_output_data)
  );
  RetimeWrapper RetimeWrapper_4 (
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_5 (
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  SingleCounter_1 SingleCounter_1 (
    .clock(SingleCounter_1_clock),
    .reset(SingleCounter_1_reset),
    .io_input_stop(SingleCounter_1_io_input_stop),
    .io_input_stride(SingleCounter_1_io_input_stride),
    .io_input_reset(SingleCounter_1_io_input_reset),
    .io_input_enable(SingleCounter_1_io_input_enable),
    .io_input_saturate(SingleCounter_1_io_input_saturate),
    .io_output_count_0(SingleCounter_1_io_output_count_0),
    .io_output_done(SingleCounter_1_io_output_done)
  );
  RetimeWrapper RetimeWrapper_6 (
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 (
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  assign _T_37 = $signed(FF_io_output_data);
  assign _T_39 = $signed(_T_37) == $signed(32'sh1);
  assign _T_40 = _T_39 & io_input_enable;
  assign _T_42 = $signed(_T_37) != $signed(32'sh1);
  assign _T_47 = _T_42 | _T_46;
  assign _T_51 = SRFF_io_output_data ? $signed(8'sh1) : $signed(8'sh2d);
  assign _T_64 = io_input_enable & io_input_stageDone_1;
  assign _T_66 = $signed(_T_63);
  assign _T_72 = $signed(_T_37) == $signed(32'sh4);
  assign _T_73 = _T_70 | _T_72;
  assign _T_91 = SingleCounter_io_output_done ? 2'h2 : 2'h1;
  assign _T_92 = {{1'd0}, _T_91};
  assign _T_96 = $signed(_T_37) < $signed(32'sh3);
  assign _T_98 = ~ io_input_stageMask_0;
  assign _T_99 = io_input_stageDone_0 | _T_98;
  assign _T_101 = ~ io_input_stageMask_1;
  assign _T_102 = io_input_stageDone_1 | _T_101;
  assign _T_104 = $signed(_T_37) - $signed(32'sh2);
  assign _T_105 = _T_104[31:0];
  assign _T_106 = $signed(_T_105);
  assign _T_107 = $unsigned(_T_106);
  assign _T_109 = 32'h1 == _T_107;
  assign _T_110 = _T_109 ? _T_102 : 1'h0;
  assign _T_111 = 32'h0 == _T_107;
  assign _T_112 = _T_111 ? _T_99 : _T_110;
  assign _T_114 = $signed(_T_37) + $signed(32'sh1);
  assign _T_115 = _T_114[31:0];
  assign _T_116 = $signed(_T_115);
  assign _T_117 = $unsigned(_T_116);
  assign _T_118 = $unsigned(_T_37);
  assign _GEN_0 = _T_112 ? _T_117 : _T_118;
  assign _T_120 = $signed(_T_37) == $signed(32'sh3);
  assign _GEN_1 = SingleCounter_1_io_output_done ? 3'h4 : 3'h2;
  assign _GEN_2 = io_input_stageDone_1 ? {{29'd0}, _GEN_1} : _T_118;
  assign _GEN_3 = _T_72 ? 32'h1 : _T_118;
  assign _GEN_4 = _T_120 ? _GEN_2 : _GEN_3;
  assign _GEN_5 = _T_96 ? _GEN_0 : _GEN_4;
  assign _GEN_6 = _T_39 ? {{29'd0}, _T_92} : _GEN_5;
  assign _GEN_8 = io_input_enable ? _GEN_6 : 32'h1;
  assign _T_144 = $signed(_T_37) == $signed(32'sh2);
  assign io_output_done = _T_72;
  assign io_output_stageEnable_0 = _T_144;
  assign io_output_stageEnable_1 = _T_120;
  assign io_output_rst_en = _T_79;
  assign SingleCounter_io_input_stop = _T_51;
  assign SingleCounter_io_input_reset = _T_47;
  assign SingleCounter_io_input_enable = _T_40;
  assign SingleCounter_clock = clock;
  assign SingleCounter_reset = reset;
  assign SRFF_io_input_set = SingleCounter_io_output_done;
  assign SRFF_io_input_reset = _T_26;
  assign SRFF_io_input_asyn_reset = _T_30;
  assign SRFF_clock = clock;
  assign SRFF_reset = reset;
  assign RetimeWrapper_io_flow = 1'h1;
  assign RetimeWrapper_io_in = reset;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_26 = RetimeWrapper_io_out;
  assign RetimeWrapper_1_io_flow = 1'h1;
  assign RetimeWrapper_1_io_in = reset;
  assign RetimeWrapper_1_clock = clock;
  assign RetimeWrapper_1_reset = reset;
  assign _T_30 = RetimeWrapper_1_io_out;
  assign FF_io_input_0_data = _GEN_8;
  assign FF_io_input_0_init = 32'h1;
  assign FF_io_input_0_enable = 1'h1;
  assign FF_io_input_0_reset = _T_36;
  assign FF_clock = clock;
  assign FF_reset = reset;
  assign RetimeWrapper_2_io_flow = 1'h1;
  assign RetimeWrapper_2_io_in = io_input_rst;
  assign RetimeWrapper_2_clock = clock;
  assign RetimeWrapper_2_reset = reset;
  assign _T_36 = RetimeWrapper_2_io_out;
  assign RetimeWrapper_3_io_flow = 1'h1;
  assign RetimeWrapper_3_io_in = io_input_rst;
  assign RetimeWrapper_3_clock = clock;
  assign RetimeWrapper_3_reset = reset;
  assign _T_46 = RetimeWrapper_3_io_out;
  assign FF_1_io_input_0_data = 32'h1;
  assign FF_1_io_input_0_init = 32'h0;
  assign FF_1_io_input_0_enable = io_input_enable;
  assign FF_1_io_input_0_reset = _T_58;
  assign FF_1_clock = clock;
  assign FF_1_reset = reset;
  assign RetimeWrapper_4_io_flow = 1'h1;
  assign RetimeWrapper_4_io_in = io_input_rst;
  assign RetimeWrapper_4_clock = clock;
  assign RetimeWrapper_4_reset = reset;
  assign _T_58 = RetimeWrapper_4_io_out;
  assign RetimeWrapper_5_io_in = FF_1_io_output_data;
  assign RetimeWrapper_5_clock = clock;
  assign RetimeWrapper_5_reset = reset;
  assign _T_63 = RetimeWrapper_5_io_out;
  assign SingleCounter_1_io_input_stop = _T_66;
  assign SingleCounter_1_io_input_stride = 32'sh0;
  assign SingleCounter_1_io_input_reset = _T_73;
  assign SingleCounter_1_io_input_enable = _T_64;
  assign SingleCounter_1_io_input_saturate = 1'h0;
  assign SingleCounter_1_clock = clock;
  assign SingleCounter_1_reset = reset;
  assign RetimeWrapper_6_io_flow = 1'h1;
  assign RetimeWrapper_6_io_in = io_input_rst;
  assign RetimeWrapper_6_clock = clock;
  assign RetimeWrapper_6_reset = reset;
  assign _T_70 = RetimeWrapper_6_io_out;
  assign RetimeWrapper_7_io_flow = 1'h1;
  assign RetimeWrapper_7_io_in = _T_39;
  assign RetimeWrapper_7_clock = clock;
  assign RetimeWrapper_7_reset = reset;
  assign _T_79 = RetimeWrapper_7_io_out;
endmodule
module SpecialAccum(
  input         clock,
  input         reset,
  input  [31:0] io_input_next,
  input         io_input_enable,
  input         io_input_reset,
  output [31:0] io_output
);
  reg [31:0] _T_10;
  reg [31:0] _RAND_0;
  wire [31:0] _T_11;
  wire [31:0] _T_13_number;
  wire [31:0] _T_15_number;
  wire [31:0] _T_17_number;
  wire [32:0] _T_19_number;
  wire [32:0] _T_21_number;
  wire [32:0] _T_23_number;
  wire [7:0] _T_27;
  wire [7:0] _T_29;
  wire [24:0] _T_31;
  wire [7:0] _T_32;
  wire  _T_33;
  wire [23:0] _T_34;
  wire [24:0] _T_35;
  wire [32:0] _T_36;
  wire [7:0] _T_40;
  wire [7:0] _T_42;
  wire [24:0] _T_44;
  wire [7:0] _T_45;
  wire  _T_46;
  wire [23:0] _T_47;
  wire [24:0] _T_48;
  wire [32:0] _T_49;
  wire [33:0] _T_50;
  wire [32:0] _T_51;
  wire [31:0] _T_53_number;
  wire [7:0] _T_63;
  wire [7:0] _T_65;
  wire [23:0] _T_67;
  wire [7:0] _T_68;
  wire [23:0] _T_70;
  wire [31:0] _T_71;
  wire [31:0] _T_72;
  assign _T_11 = io_input_reset ? 32'h0 : _T_10;
  assign _T_32 = _T_15_number[7:0];
  assign _T_33 = _T_15_number[31];
  assign _T_34 = _T_15_number[31:8];
  assign _T_35 = {_T_33,_T_34};
  assign _T_36 = {_T_31,_T_29};
  assign _T_45 = _T_13_number[7:0];
  assign _T_46 = _T_13_number[31];
  assign _T_47 = _T_13_number[31:8];
  assign _T_48 = {_T_46,_T_47};
  assign _T_49 = {_T_44,_T_42};
  assign _T_50 = _T_21_number + _T_23_number;
  assign _T_51 = _T_50[32:0];
  assign _T_68 = _T_19_number[7:0];
  assign _T_70 = _T_19_number[31:8];
  assign _T_71 = {_T_67,_T_65};
  assign _T_72 = io_input_enable ? _T_53_number : _T_17_number;
  assign io_output = _T_11;
  assign _T_13_number = io_input_next;
  assign _T_15_number = _T_10;
  assign _T_17_number = _T_11;
  assign _T_19_number = _T_51;
  assign _T_21_number = _T_36;
  assign _T_23_number = _T_49;
  assign _T_27 = _T_32;
  assign _T_29 = _T_27;
  assign _T_31 = _T_35;
  assign _T_40 = _T_45;
  assign _T_42 = _T_40;
  assign _T_44 = _T_48;
  assign _T_53_number = _T_71;
  assign _T_63 = _T_68;
  assign _T_65 = _T_63;
  assign _T_67 = _T_70;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_10 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_10 <= 32'h0;
    end else begin
      if (io_input_enable) begin
        _T_10 <= _T_53_number;
      end else begin
        _T_10 <= _T_17_number;
      end
    end
  end
endmodule
module SingleCounter_2(
  input         clock,
  input         reset,
  input  [31:0] io_input_stop,
  input         io_input_reset,
  input         io_input_enable,
  output [31:0] io_output_count_0,
  output [31:0] io_output_count_1
);
  wire  FF_clock;
  wire  FF_reset;
  wire [31:0] FF_io_input_0_data;
  wire [31:0] FF_io_input_0_init;
  wire  FF_io_input_0_enable;
  wire  FF_io_input_0_reset;
  wire [31:0] FF_io_output_data;
  wire  FF_1_clock;
  wire  FF_1_reset;
  wire [31:0] FF_1_io_input_0_data;
  wire [31:0] FF_1_io_input_0_init;
  wire  FF_1_io_input_0_enable;
  wire  FF_1_io_input_0_reset;
  wire [31:0] FF_1_io_output_data;
  wire [31:0] _T_24;
  wire [31:0] _T_25;
  wire [32:0] _T_27;
  wire [31:0] _T_28;
  wire [31:0] _T_29;
  wire [32:0] _T_30;
  wire [31:0] _T_31;
  wire [31:0] _T_32;
  wire  _T_35;
  wire [31:0] _T_48;
  wire [31:0] _T_49;
  wire [31:0] _T_50;
  wire [31:0] _T_55;
  wire [31:0] _T_56;
  wire [31:0] _T_57;
  FF_1 FF (
    .clock(FF_clock),
    .reset(FF_reset),
    .io_input_0_data(FF_io_input_0_data),
    .io_input_0_init(FF_io_input_0_init),
    .io_input_0_enable(FF_io_input_0_enable),
    .io_input_0_reset(FF_io_input_0_reset),
    .io_output_data(FF_io_output_data)
  );
  FF_1 FF_1 (
    .clock(FF_1_clock),
    .reset(FF_1_reset),
    .io_input_0_data(FF_1_io_input_0_data),
    .io_input_0_init(FF_1_io_input_0_init),
    .io_input_0_enable(FF_1_io_input_0_enable),
    .io_input_0_reset(FF_1_io_input_0_reset),
    .io_output_data(FF_1_io_output_data)
  );
  assign _T_24 = $signed(FF_io_output_data);
  assign _T_25 = $signed(FF_1_io_output_data);
  assign _T_27 = $signed(_T_24) + $signed(32'sh80);
  assign _T_28 = _T_27[31:0];
  assign _T_29 = $signed(_T_28);
  assign _T_30 = $signed(_T_25) + $signed(32'sh80);
  assign _T_31 = _T_30[31:0];
  assign _T_32 = $signed(_T_31);
  assign _T_35 = $signed(_T_29) >= $signed(io_input_stop);
  assign _T_48 = $unsigned(_T_29);
  assign _T_49 = _T_35 ? 32'h0 : _T_48;
  assign _T_50 = io_input_reset ? 32'h0 : _T_49;
  assign _T_55 = $unsigned(_T_32);
  assign _T_56 = _T_35 ? 32'h40 : _T_55;
  assign _T_57 = io_input_reset ? 32'h40 : _T_56;
  assign io_output_count_0 = _T_24;
  assign io_output_count_1 = _T_25;
  assign FF_io_input_0_data = _T_50;
  assign FF_io_input_0_init = 32'h0;
  assign FF_io_input_0_enable = io_input_enable;
  assign FF_io_input_0_reset = io_input_reset;
  assign FF_clock = clock;
  assign FF_reset = reset;
  assign FF_1_io_input_0_data = _T_57;
  assign FF_1_io_input_0_init = 32'h40;
  assign FF_1_io_input_0_enable = io_input_enable;
  assign FF_1_io_input_0_reset = io_input_reset;
  assign FF_1_clock = clock;
  assign FF_1_reset = reset;
endmodule
module Counter(
  input         clock,
  input         reset,
  input  [31:0] io_input_stops_0,
  input         io_input_reset,
  input         io_input_enable,
  output [31:0] io_output_counts_1,
  output [31:0] io_output_counts_0
);
  wire  ctrs_0_clock;
  wire  ctrs_0_reset;
  wire [31:0] ctrs_0_io_input_stop;
  wire  ctrs_0_io_input_reset;
  wire  ctrs_0_io_input_enable;
  wire [31:0] ctrs_0_io_output_count_0;
  wire [31:0] ctrs_0_io_output_count_1;
  SingleCounter_2 ctrs_0 (
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_input_stop(ctrs_0_io_input_stop),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_count_1(ctrs_0_io_output_count_1)
  );
  assign io_output_counts_1 = ctrs_0_io_output_count_1;
  assign io_output_counts_0 = ctrs_0_io_output_count_0;
  assign ctrs_0_io_input_stop = io_input_stops_0;
  assign ctrs_0_io_input_reset = io_input_reset;
  assign ctrs_0_io_input_enable = io_input_enable;
  assign ctrs_0_clock = clock;
  assign ctrs_0_reset = reset;
endmodule
module FF_11(
  input        clock,
  input        reset,
  input  [2:0] io_input_0_data,
  input        io_input_0_enable,
  input        io_input_0_reset,
  output [2:0] io_output_data
);
  reg [2:0] ff;
  reg [31:0] _RAND_0;
  wire [2:0] _T_7;
  wire [2:0] _T_8;
  wire [2:0] _T_9;
  assign _T_7 = io_input_0_enable ? io_input_0_data : ff;
  assign _T_8 = io_input_0_reset ? 3'h0 : _T_7;
  assign _T_9 = io_input_0_reset ? 3'h0 : ff;
  assign io_output_data = _T_9;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  ff = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 3'h0;
    end else begin
      if (io_input_0_reset) begin
        ff <= 3'h0;
      end else begin
        if (io_input_0_enable) begin
          ff <= io_input_0_data;
        end
      end
    end
  end
endmodule
module Metapipe(
  input         clock,
  input         reset,
  input         io_input_enable,
  input  [31:0] io_input_numIter,
  input         io_input_stageDone_0,
  input         io_input_stageDone_1,
  input         io_input_stageDone_2,
  input         io_input_stageDone_3,
  input         io_input_stageDone_4,
  input         io_input_rst,
  output        io_output_done,
  output        io_output_stageEnable_0,
  output        io_output_stageEnable_1,
  output        io_output_stageEnable_2,
  output        io_output_stageEnable_3,
  output        io_output_stageEnable_4,
  output        io_output_rst_en,
  output        io_output_ctr_inc
);
  wire  deadState_clock;
  wire  deadState_reset;
  wire  deadState_io_input_set;
  wire  deadState_io_input_reset;
  wire  deadState_io_input_asyn_reset;
  wire  deadState_io_output_data;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire  RetimeWrapper_io_flow;
  wire  RetimeWrapper_io_in;
  wire  RetimeWrapper_io_out;
  wire  _T_24;
  wire  rstCtr_clock;
  wire  rstCtr_reset;
  wire [7:0] rstCtr_io_input_stop;
  wire  rstCtr_io_input_reset;
  wire  rstCtr_io_input_enable;
  wire  rstCtr_io_output_done;
  wire  firstIterComplete_clock;
  wire  firstIterComplete_reset;
  wire  firstIterComplete_io_input_set;
  wire  firstIterComplete_io_input_reset;
  wire  firstIterComplete_io_input_asyn_reset;
  wire  firstIterComplete_io_output_data;
  wire  RetimeWrapper_1_clock;
  wire  RetimeWrapper_1_reset;
  wire  RetimeWrapper_1_io_flow;
  wire  RetimeWrapper_1_io_in;
  wire  RetimeWrapper_1_io_out;
  wire  _T_28;
  wire  RetimeWrapper_2_clock;
  wire  RetimeWrapper_2_reset;
  wire  RetimeWrapper_2_io_flow;
  wire  RetimeWrapper_2_io_in;
  wire  RetimeWrapper_2_io_out;
  wire  _T_32;
  wire  stateFF_clock;
  wire  stateFF_reset;
  wire [31:0] stateFF_io_input_0_data;
  wire [31:0] stateFF_io_input_0_init;
  wire  stateFF_io_input_0_enable;
  wire  stateFF_io_input_0_reset;
  wire [31:0] stateFF_io_output_data;
  wire  RetimeWrapper_3_clock;
  wire  RetimeWrapper_3_reset;
  wire  RetimeWrapper_3_io_flow;
  wire  RetimeWrapper_3_io_in;
  wire  RetimeWrapper_3_io_out;
  wire  _T_38;
  wire  _T_40;
  wire  _T_41;
  wire  _T_43;
  wire  RetimeWrapper_4_clock;
  wire  RetimeWrapper_4_reset;
  wire  RetimeWrapper_4_io_flow;
  wire  RetimeWrapper_4_io_in;
  wire  RetimeWrapper_4_io_out;
  wire  _T_47;
  wire  _T_48;
  wire  maxFF_clock;
  wire  maxFF_reset;
  wire [31:0] maxFF_io_input_0_data;
  wire [31:0] maxFF_io_input_0_init;
  wire  maxFF_io_input_0_enable;
  wire  maxFF_io_input_0_reset;
  wire [31:0] maxFF_io_output_data;
  wire  RetimeWrapper_5_clock;
  wire  RetimeWrapper_5_reset;
  wire  RetimeWrapper_5_io_flow;
  wire  RetimeWrapper_5_io_in;
  wire  RetimeWrapper_5_io_out;
  wire  _T_63;
  wire  RetimeWrapper_6_clock;
  wire  RetimeWrapper_6_reset;
  wire [31:0] RetimeWrapper_6_io_in;
  wire [31:0] RetimeWrapper_6_io_out;
  wire [31:0] max;
  wire  doneClear;
  wire  doneFF_0_clock;
  wire  doneFF_0_reset;
  wire  doneFF_0_io_input_set;
  wire  doneFF_0_io_input_reset;
  wire  doneFF_0_io_input_asyn_reset;
  wire  doneFF_0_io_output_data;
  wire  RetimeWrapper_7_clock;
  wire  RetimeWrapper_7_reset;
  wire  RetimeWrapper_7_io_flow;
  wire  RetimeWrapper_7_io_in;
  wire  RetimeWrapper_7_io_out;
  wire  _T_71;
  wire  doneFF_1_clock;
  wire  doneFF_1_reset;
  wire  doneFF_1_io_input_set;
  wire  doneFF_1_io_input_reset;
  wire  doneFF_1_io_input_asyn_reset;
  wire  doneFF_1_io_output_data;
  wire  RetimeWrapper_8_clock;
  wire  RetimeWrapper_8_reset;
  wire  RetimeWrapper_8_io_flow;
  wire  RetimeWrapper_8_io_in;
  wire  RetimeWrapper_8_io_out;
  wire  _T_75;
  wire  doneFF_2_clock;
  wire  doneFF_2_reset;
  wire  doneFF_2_io_input_set;
  wire  doneFF_2_io_input_reset;
  wire  doneFF_2_io_input_asyn_reset;
  wire  doneFF_2_io_output_data;
  wire  RetimeWrapper_9_clock;
  wire  RetimeWrapper_9_reset;
  wire  RetimeWrapper_9_io_flow;
  wire  RetimeWrapper_9_io_in;
  wire  RetimeWrapper_9_io_out;
  wire  _T_79;
  wire  doneFF_3_clock;
  wire  doneFF_3_reset;
  wire  doneFF_3_io_input_set;
  wire  doneFF_3_io_input_reset;
  wire  doneFF_3_io_input_asyn_reset;
  wire  doneFF_3_io_output_data;
  wire  RetimeWrapper_10_clock;
  wire  RetimeWrapper_10_reset;
  wire  RetimeWrapper_10_io_flow;
  wire  RetimeWrapper_10_io_in;
  wire  RetimeWrapper_10_io_out;
  wire  _T_83;
  wire  doneFF_4_clock;
  wire  doneFF_4_reset;
  wire  doneFF_4_io_input_set;
  wire  doneFF_4_io_input_reset;
  wire  doneFF_4_io_input_asyn_reset;
  wire  doneFF_4_io_output_data;
  wire  RetimeWrapper_11_clock;
  wire  RetimeWrapper_11_reset;
  wire  RetimeWrapper_11_io_flow;
  wire  RetimeWrapper_11_io_in;
  wire  RetimeWrapper_11_io_out;
  wire  _T_87;
  wire  ctr_clock;
  wire  ctr_reset;
  wire [31:0] ctr_io_input_stop;
  wire [31:0] ctr_io_input_stride;
  wire  ctr_io_input_reset;
  wire  ctr_io_input_enable;
  wire  ctr_io_input_saturate;
  wire [31:0] ctr_io_output_count_0;
  wire  ctr_io_output_done;
  wire [31:0] _T_89;
  wire  _T_91;
  wire  _T_92;
  wire  RetimeWrapper_12_clock;
  wire  RetimeWrapper_12_reset;
  wire  RetimeWrapper_12_io_flow;
  wire  RetimeWrapper_12_io_in;
  wire  RetimeWrapper_12_io_out;
  wire  _T_96;
  wire  RetimeWrapper_13_clock;
  wire  RetimeWrapper_13_reset;
  wire  RetimeWrapper_13_io_flow;
  wire  RetimeWrapper_13_io_in;
  wire  RetimeWrapper_13_io_out;
  wire  _T_102;
  wire  cycsSinceDone_clock;
  wire  cycsSinceDone_reset;
  wire [2:0] cycsSinceDone_io_input_0_data;
  wire  cycsSinceDone_io_input_0_enable;
  wire  cycsSinceDone_io_input_0_reset;
  wire [2:0] cycsSinceDone_io_output_data;
  wire  _T_111;
  wire [3:0] _T_115;
  wire [1:0] _T_119;
  wire [3:0] _T_120;
  wire  _T_128;
  wire  _T_131;
  wire  _T_133;
  wire  _T_134;
  wire  _T_136;
  wire  _T_137;
  wire  _T_144;
  wire  _T_147;
  wire  _T_149;
  wire  _T_151;
  wire  _T_152;
  wire  _T_154;
  wire  _T_156;
  wire  _T_157;
  wire  _T_159;
  wire  _T_161;
  wire  _T_162;
  wire  _T_164;
  wire [2:0] _T_170;
  wire [3:0] _T_171;
  wire [2:0] _T_172;
  wire  _T_174;
  wire [3:0] _T_178;
  wire [2:0] _T_179;
  wire [32:0] _T_181;
  wire [31:0] _T_182;
  wire [31:0] _T_183;
  wire  _T_185;
  wire  _GEN_1;
  wire [31:0] _GEN_3;
  wire  _T_191;
  wire  _T_200;
  wire  _T_203;
  wire  _T_206;
  wire [2:0] _T_241;
  wire [3:0] _T_242;
  wire [2:0] _T_243;
  wire [3:0] _T_244;
  wire [2:0] _T_245;
  wire  _T_247;
  wire [2:0] _GEN_11;
  wire  _GEN_12;
  wire [31:0] _GEN_14;
  wire  _GEN_15;
  wire  _GEN_16;
  wire  _GEN_18;
  wire [2:0] _GEN_19;
  wire  _GEN_20;
  wire [31:0] _GEN_22;
  wire  _T_264;
  wire  _T_281;
  wire  _T_284;
  wire  _T_287;
  wire [2:0] _T_324;
  wire [3:0] _T_327;
  wire [2:0] _T_328;
  wire [3:0] _T_329;
  wire [2:0] _T_330;
  wire  _T_332;
  wire [2:0] _GEN_23;
  wire  _GEN_24;
  wire [31:0] _GEN_26;
  wire  _GEN_27;
  wire  _GEN_28;
  wire  _GEN_29;
  wire  _GEN_31;
  wire [2:0] _GEN_32;
  wire  _GEN_33;
  wire [31:0] _GEN_35;
  wire  _T_349;
  wire  _T_374;
  wire  _T_377;
  wire  _T_380;
  wire [2:0] _T_419;
  wire [3:0] _T_424;
  wire [2:0] _T_425;
  wire [3:0] _T_426;
  wire [2:0] _T_427;
  wire  _T_429;
  wire  _T_434;
  wire  _T_440;
  wire  _T_441;
  wire [3:0] _T_445;
  wire [2:0] _T_446;
  wire [31:0] _GEN_144;
  wire [32:0] _T_447;
  wire [31:0] _T_448;
  wire [31:0] _T_450;
  wire [31:0] _GEN_37;
  wire  _GEN_39;
  wire  _GEN_40;
  wire  _GEN_41;
  wire  _GEN_42;
  wire  _GEN_44;
  wire  _GEN_45;
  wire [31:0] _GEN_46;
  wire  _T_455;
  wire  _T_464;
  wire  _T_477;
  wire  _T_478;
  wire  _T_479;
  wire  _T_480;
  wire  RetimeWrapper_14_clock;
  wire  RetimeWrapper_14_reset;
  wire [31:0] RetimeWrapper_14_io_in;
  wire [31:0] RetimeWrapper_14_io_out;
  wire [31:0] _T_484;
  wire [31:0] _T_487;
  wire [31:0] _T_488;
  wire [32:0] _T_491;
  wire [31:0] _T_492;
  wire [31:0] _T_493;
  wire  _T_494;
  wire [31:0] _GEN_48;
  wire [31:0] _GEN_50;
  wire  _GEN_51;
  wire  _T_502;
  wire  _T_525;
  wire  _T_526;
  wire  _T_527;
  wire [31:0] _GEN_52;
  wire  _T_534;
  wire  _T_553;
  wire  _T_554;
  wire [31:0] _GEN_62;
  wire  _GEN_64;
  wire  _GEN_65;
  wire  _GEN_66;
  wire  _GEN_68;
  wire  _GEN_69;
  wire [31:0] _GEN_70;
  wire  _T_561;
  wire  _T_579;
  wire [31:0] _GEN_72;
  wire  _GEN_74;
  wire  _GEN_75;
  wire  _GEN_77;
  wire  _GEN_78;
  wire  _GEN_79;
  wire [31:0] _GEN_80;
  wire  _T_586;
  wire [31:0] _GEN_82;
  wire  _GEN_84;
  wire  _GEN_86;
  wire  _GEN_87;
  wire  _GEN_88;
  wire  _GEN_89;
  wire [31:0] _GEN_90;
  wire [31:0] _GEN_94;
  wire  _GEN_96;
  wire  _GEN_97;
  wire  _GEN_98;
  wire  _GEN_99;
  wire  _GEN_101;
  wire [31:0] _GEN_102;
  wire  _GEN_104;
  wire  _GEN_105;
  wire  _GEN_106;
  wire  _GEN_107;
  wire  _GEN_108;
  wire  _GEN_110;
  wire [31:0] _GEN_111;
  wire  _GEN_112;
  wire  _GEN_113;
  wire  _GEN_114;
  wire  _GEN_115;
  wire  _GEN_116;
  wire  _GEN_117;
  wire  _GEN_118;
  wire  _GEN_120;
  wire  _GEN_121;
  wire [31:0] _GEN_122;
  wire  _GEN_123;
  wire [31:0] _GEN_124;
  wire  _GEN_125;
  wire  _GEN_126;
  wire  _GEN_127;
  wire  _GEN_128;
  wire  _GEN_129;
  wire  _GEN_130;
  wire  _GEN_133;
  wire  _GEN_134;
  wire [31:0] _GEN_135;
  wire  _GEN_136;
  wire  _GEN_137;
  wire  _GEN_138;
  wire  _GEN_139;
  wire  _GEN_140;
  wire  _GEN_141;
  wire  _GEN_143;
  wire  _T_634;
  reg  _T_637;
  reg [31:0] _RAND_0;
  wire  _T_643;
  SRFF deadState (
    .clock(deadState_clock),
    .reset(deadState_reset),
    .io_input_set(deadState_io_input_set),
    .io_input_reset(deadState_io_input_reset),
    .io_input_asyn_reset(deadState_io_input_asyn_reset),
    .io_output_data(deadState_io_output_data)
  );
  RetimeWrapper RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  SingleCounter rstCtr (
    .clock(rstCtr_clock),
    .reset(rstCtr_reset),
    .io_input_stop(rstCtr_io_input_stop),
    .io_input_reset(rstCtr_io_input_reset),
    .io_input_enable(rstCtr_io_input_enable),
    .io_output_done(rstCtr_io_output_done)
  );
  SRFF firstIterComplete (
    .clock(firstIterComplete_clock),
    .reset(firstIterComplete_reset),
    .io_input_set(firstIterComplete_io_input_set),
    .io_input_reset(firstIterComplete_io_input_reset),
    .io_input_asyn_reset(firstIterComplete_io_input_asyn_reset),
    .io_output_data(firstIterComplete_io_output_data)
  );
  RetimeWrapper RetimeWrapper_1 (
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 (
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  FF_1 stateFF (
    .clock(stateFF_clock),
    .reset(stateFF_reset),
    .io_input_0_data(stateFF_io_input_0_data),
    .io_input_0_init(stateFF_io_input_0_init),
    .io_input_0_enable(stateFF_io_input_0_enable),
    .io_input_0_reset(stateFF_io_input_0_reset),
    .io_output_data(stateFF_io_output_data)
  );
  RetimeWrapper RetimeWrapper_3 (
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 (
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  FF_1 maxFF (
    .clock(maxFF_clock),
    .reset(maxFF_reset),
    .io_input_0_data(maxFF_io_input_0_data),
    .io_input_0_init(maxFF_io_input_0_init),
    .io_input_0_enable(maxFF_io_input_0_enable),
    .io_input_0_reset(maxFF_io_input_0_reset),
    .io_output_data(maxFF_io_output_data)
  );
  RetimeWrapper RetimeWrapper_5 (
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_6 (
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  SRFF doneFF_0 (
    .clock(doneFF_0_clock),
    .reset(doneFF_0_reset),
    .io_input_set(doneFF_0_io_input_set),
    .io_input_reset(doneFF_0_io_input_reset),
    .io_input_asyn_reset(doneFF_0_io_input_asyn_reset),
    .io_output_data(doneFF_0_io_output_data)
  );
  RetimeWrapper RetimeWrapper_7 (
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  SRFF doneFF_1 (
    .clock(doneFF_1_clock),
    .reset(doneFF_1_reset),
    .io_input_set(doneFF_1_io_input_set),
    .io_input_reset(doneFF_1_io_input_reset),
    .io_input_asyn_reset(doneFF_1_io_input_asyn_reset),
    .io_output_data(doneFF_1_io_output_data)
  );
  RetimeWrapper RetimeWrapper_8 (
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  SRFF doneFF_2 (
    .clock(doneFF_2_clock),
    .reset(doneFF_2_reset),
    .io_input_set(doneFF_2_io_input_set),
    .io_input_reset(doneFF_2_io_input_reset),
    .io_input_asyn_reset(doneFF_2_io_input_asyn_reset),
    .io_output_data(doneFF_2_io_output_data)
  );
  RetimeWrapper RetimeWrapper_9 (
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  SRFF doneFF_3 (
    .clock(doneFF_3_clock),
    .reset(doneFF_3_reset),
    .io_input_set(doneFF_3_io_input_set),
    .io_input_reset(doneFF_3_io_input_reset),
    .io_input_asyn_reset(doneFF_3_io_input_asyn_reset),
    .io_output_data(doneFF_3_io_output_data)
  );
  RetimeWrapper RetimeWrapper_10 (
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  SRFF doneFF_4 (
    .clock(doneFF_4_clock),
    .reset(doneFF_4_reset),
    .io_input_set(doneFF_4_io_input_set),
    .io_input_reset(doneFF_4_io_input_reset),
    .io_input_asyn_reset(doneFF_4_io_input_asyn_reset),
    .io_output_data(doneFF_4_io_output_data)
  );
  RetimeWrapper RetimeWrapper_11 (
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  SingleCounter_1 ctr (
    .clock(ctr_clock),
    .reset(ctr_reset),
    .io_input_stop(ctr_io_input_stop),
    .io_input_stride(ctr_io_input_stride),
    .io_input_reset(ctr_io_input_reset),
    .io_input_enable(ctr_io_input_enable),
    .io_input_saturate(ctr_io_input_saturate),
    .io_output_count_0(ctr_io_output_count_0),
    .io_output_done(ctr_io_output_done)
  );
  RetimeWrapper RetimeWrapper_12 (
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper RetimeWrapper_13 (
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  FF_11 cycsSinceDone (
    .clock(cycsSinceDone_clock),
    .reset(cycsSinceDone_reset),
    .io_input_0_data(cycsSinceDone_io_input_0_data),
    .io_input_0_enable(cycsSinceDone_io_input_0_enable),
    .io_input_0_reset(cycsSinceDone_io_input_0_reset),
    .io_output_data(cycsSinceDone_io_output_data)
  );
  RetimeWrapper_6 RetimeWrapper_14 (
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  assign _T_40 = stateFF_io_output_data == 32'h1;
  assign _T_41 = _T_40 & io_input_enable;
  assign _T_43 = stateFF_io_output_data != 32'h1;
  assign _T_48 = _T_43 | _T_47;
  assign _T_89 = $signed(max);
  assign _T_91 = stateFF_io_output_data == 32'hb;
  assign _T_92 = io_input_rst | _T_91;
  assign _T_111 = io_input_numIter == 32'h0;
  assign _T_115 = rstCtr_io_output_done ? 4'hb : 4'h1;
  assign _T_119 = rstCtr_io_output_done ? 2'h2 : 2'h1;
  assign _T_120 = _T_111 ? _T_115 : {{2'd0}, _T_119};
  assign _T_128 = stateFF_io_output_data < 32'h6;
  assign _T_131 = ~ doneFF_0_io_output_data;
  assign _T_133 = 3'h0 >= cycsSinceDone_io_output_data;
  assign _T_134 = _T_131 & _T_133;
  assign _T_136 = io_input_numIter != 32'h0;
  assign _T_137 = _T_134 & _T_136;
  assign _T_144 = doneFF_0_io_output_data;
  assign _T_147 = _T_144 & _T_133;
  assign _T_149 = doneFF_1_io_output_data;
  assign _T_151 = 3'h1 >= cycsSinceDone_io_output_data;
  assign _T_152 = _T_149 & _T_151;
  assign _T_154 = doneFF_2_io_output_data;
  assign _T_156 = 3'h2 >= cycsSinceDone_io_output_data;
  assign _T_157 = _T_154 & _T_156;
  assign _T_159 = doneFF_3_io_output_data;
  assign _T_161 = 3'h3 >= cycsSinceDone_io_output_data;
  assign _T_162 = _T_159 & _T_161;
  assign _T_164 = doneFF_4_io_output_data;
  assign _T_170 = _T_147 ? 3'h1 : 3'h0;
  assign _T_171 = _T_170 + cycsSinceDone_io_output_data;
  assign _T_172 = _T_171[2:0];
  assign _T_174 = _T_172 == 3'h1;
  assign _T_178 = cycsSinceDone_io_output_data + 3'h1;
  assign _T_179 = _T_178[2:0];
  assign _T_181 = $signed(ctr_io_output_count_0) + $signed(32'sh1);
  assign _T_182 = _T_181[31:0];
  assign _T_183 = $signed(_T_182);
  assign _T_185 = $signed(_T_183) == $signed(_T_89);
  assign _GEN_1 = _T_174 ? _T_185 : 1'h0;
  assign _GEN_3 = _T_174 ? 32'h3 : stateFF_io_output_data;
  assign _T_191 = stateFF_io_output_data == 32'h3;
  assign _T_200 = ~ doneFF_1_io_output_data;
  assign _T_203 = _T_200 & _T_151;
  assign _T_206 = _T_203 & _T_136;
  assign _T_241 = _T_152 ? 3'h1 : 3'h0;
  assign _T_242 = _T_170 + _T_241;
  assign _T_243 = _T_242[2:0];
  assign _T_244 = _T_243 + cycsSinceDone_io_output_data;
  assign _T_245 = _T_244[2:0];
  assign _T_247 = _T_245 == 3'h2;
  assign _GEN_11 = _T_247 ? _T_179 : _T_179;
  assign _GEN_12 = _T_247 ? _T_185 : 1'h0;
  assign _GEN_14 = _T_247 ? 32'h4 : stateFF_io_output_data;
  assign _GEN_15 = _T_191 ? _T_137 : _T_137;
  assign _GEN_16 = _T_191 ? _T_206 : 1'h0;
  assign _GEN_18 = _T_191 ? _T_247 : _T_174;
  assign _GEN_19 = _T_191 ? _GEN_11 : _T_179;
  assign _GEN_20 = _T_191 ? _GEN_12 : _GEN_1;
  assign _GEN_22 = _T_191 ? _GEN_14 : _GEN_3;
  assign _T_264 = stateFF_io_output_data == 32'h4;
  assign _T_281 = ~ doneFF_2_io_output_data;
  assign _T_284 = _T_281 & _T_156;
  assign _T_287 = _T_284 & _T_136;
  assign _T_324 = _T_157 ? 3'h1 : 3'h0;
  assign _T_327 = _T_243 + _T_324;
  assign _T_328 = _T_327[2:0];
  assign _T_329 = _T_328 + cycsSinceDone_io_output_data;
  assign _T_330 = _T_329[2:0];
  assign _T_332 = _T_330 == 3'h3;
  assign _GEN_23 = _T_332 ? _T_179 : _GEN_19;
  assign _GEN_24 = _T_332 ? _T_185 : 1'h0;
  assign _GEN_26 = _T_332 ? 32'h5 : stateFF_io_output_data;
  assign _GEN_27 = _T_264 ? _T_137 : _GEN_15;
  assign _GEN_28 = _T_264 ? _T_206 : _GEN_16;
  assign _GEN_29 = _T_264 ? _T_287 : 1'h0;
  assign _GEN_31 = _T_264 ? _T_332 : _GEN_18;
  assign _GEN_32 = _T_264 ? _GEN_23 : _GEN_19;
  assign _GEN_33 = _T_264 ? _GEN_24 : _GEN_20;
  assign _GEN_35 = _T_264 ? _GEN_26 : _GEN_22;
  assign _T_349 = stateFF_io_output_data == 32'h5;
  assign _T_374 = ~ doneFF_3_io_output_data;
  assign _T_377 = _T_374 & _T_161;
  assign _T_380 = _T_377 & _T_136;
  assign _T_419 = _T_162 ? 3'h1 : 3'h0;
  assign _T_424 = _T_328 + _T_419;
  assign _T_425 = _T_424[2:0];
  assign _T_426 = _T_425 + cycsSinceDone_io_output_data;
  assign _T_427 = _T_426[2:0];
  assign _T_429 = _T_427 == 3'h4;
  assign _T_434 = cycsSinceDone_io_output_data == 3'h0;
  assign _T_440 = $signed(_T_183) < $signed(_T_89);
  assign _T_441 = _T_434 & _T_440;
  assign _T_445 = cycsSinceDone_io_output_data + 3'h2;
  assign _T_446 = _T_445[2:0];
  assign _GEN_144 = {{29'd0}, _T_446};
  assign _T_447 = _GEN_144 + stateFF_io_output_data;
  assign _T_448 = _T_447[31:0];
  assign _T_450 = _T_441 ? 32'h6 : _T_448;
  assign _GEN_37 = _T_429 ? _T_450 : stateFF_io_output_data;
  assign _GEN_39 = _T_349 ? _T_137 : _GEN_27;
  assign _GEN_40 = _T_349 ? _T_206 : _GEN_28;
  assign _GEN_41 = _T_349 ? _T_287 : _GEN_29;
  assign _GEN_42 = _T_349 ? _T_380 : 1'h0;
  assign _GEN_44 = _T_349 ? _T_429 : _GEN_31;
  assign _GEN_45 = _T_349 ? 1'h0 : _GEN_33;
  assign _GEN_46 = _T_349 ? _GEN_37 : _GEN_35;
  assign _T_455 = stateFF_io_output_data == 32'h6;
  assign _T_464 = ~ doneFF_4_io_output_data;
  assign _T_477 = _T_144 & _T_149;
  assign _T_478 = _T_477 & _T_154;
  assign _T_479 = _T_478 & _T_159;
  assign _T_480 = _T_479 & _T_164;
  assign _T_484 = $unsigned(ctr_io_output_count_0);
  assign _T_488 = $signed(RetimeWrapper_14_io_out);
  assign _T_491 = $signed(_T_89) - $signed(32'sh1);
  assign _T_492 = _T_491[31:0];
  assign _T_493 = $signed(_T_492);
  assign _T_494 = $signed(_T_487) == $signed(_T_493);
  assign _GEN_48 = _T_494 ? 32'h7 : stateFF_io_output_data;
  assign _GEN_50 = _T_480 ? _GEN_48 : stateFF_io_output_data;
  assign _GEN_51 = _T_480 ? _T_494 : 1'h0;
  assign _T_502 = stateFF_io_output_data < 32'hb;
  assign _T_525 = _T_149 & _T_154;
  assign _T_526 = _T_525 & _T_159;
  assign _T_527 = _T_526 & _T_164;
  assign _GEN_52 = _T_527 ? 32'h8 : stateFF_io_output_data;
  assign _T_534 = stateFF_io_output_data == 32'h8;
  assign _T_553 = _T_154 & _T_159;
  assign _T_554 = _T_553 & _T_164;
  assign _GEN_62 = _T_554 ? 32'h9 : stateFF_io_output_data;
  assign _GEN_64 = _T_534 ? _T_281 : _T_281;
  assign _GEN_65 = _T_534 ? _T_374 : _T_374;
  assign _GEN_66 = _T_534 ? _T_464 : _T_464;
  assign _GEN_68 = _T_534 ? 1'h0 : _T_200;
  assign _GEN_69 = _T_534 ? _T_554 : _T_527;
  assign _GEN_70 = _T_534 ? _GEN_62 : _GEN_52;
  assign _T_561 = stateFF_io_output_data == 32'h9;
  assign _T_579 = _T_159 & _T_164;
  assign _GEN_72 = _T_579 ? 32'ha : stateFF_io_output_data;
  assign _GEN_74 = _T_561 ? _T_374 : _GEN_65;
  assign _GEN_75 = _T_561 ? _T_464 : _GEN_66;
  assign _GEN_77 = _T_561 ? 1'h0 : _GEN_68;
  assign _GEN_78 = _T_561 ? 1'h0 : _GEN_64;
  assign _GEN_79 = _T_561 ? _T_579 : _GEN_69;
  assign _GEN_80 = _T_561 ? _GEN_72 : _GEN_70;
  assign _T_586 = stateFF_io_output_data == 32'ha;
  assign _GEN_82 = _T_164 ? 32'hb : stateFF_io_output_data;
  assign _GEN_84 = _T_586 ? _T_464 : _GEN_75;
  assign _GEN_86 = _T_586 ? 1'h0 : _GEN_77;
  assign _GEN_87 = _T_586 ? 1'h0 : _GEN_78;
  assign _GEN_88 = _T_586 ? 1'h0 : _GEN_74;
  assign _GEN_89 = _T_586 ? _T_164 : _GEN_79;
  assign _GEN_90 = _T_586 ? _GEN_82 : _GEN_80;
  assign _GEN_94 = _T_91 ? 32'h1 : stateFF_io_output_data;
  assign _GEN_96 = _T_502 ? _GEN_86 : 1'h0;
  assign _GEN_97 = _T_502 ? _GEN_87 : 1'h0;
  assign _GEN_98 = _T_502 ? _GEN_88 : 1'h0;
  assign _GEN_99 = _T_502 ? _GEN_84 : 1'h0;
  assign _GEN_101 = _T_502 ? _GEN_89 : 1'h0;
  assign _GEN_102 = _T_502 ? _GEN_90 : _GEN_94;
  assign _GEN_104 = _T_455 ? _T_131 : 1'h0;
  assign _GEN_105 = _T_455 ? _T_200 : _GEN_96;
  assign _GEN_106 = _T_455 ? _T_281 : _GEN_97;
  assign _GEN_107 = _T_455 ? _T_374 : _GEN_98;
  assign _GEN_108 = _T_455 ? _T_464 : _GEN_99;
  assign _GEN_110 = _T_455 ? _T_480 : _GEN_101;
  assign _GEN_111 = _T_455 ? _GEN_50 : _GEN_102;
  assign _GEN_112 = _T_455 ? _GEN_51 : _GEN_101;
  assign _GEN_113 = _T_128 ? _GEN_39 : _GEN_104;
  assign _GEN_114 = _T_128 ? _GEN_40 : _GEN_105;
  assign _GEN_115 = _T_128 ? _GEN_41 : _GEN_106;
  assign _GEN_116 = _T_128 ? _GEN_42 : _GEN_107;
  assign _GEN_117 = _T_128 ? 1'h0 : _GEN_108;
  assign _GEN_118 = _T_128 ? _GEN_44 : _GEN_110;
  assign _GEN_120 = _T_128 ? _GEN_45 : 1'h0;
  assign _GEN_121 = _T_128 ? _GEN_44 : _GEN_112;
  assign _GEN_122 = _T_128 ? _GEN_46 : _GEN_111;
  assign _GEN_123 = _T_40 ? 1'h0 : _GEN_118;
  assign _GEN_124 = _T_40 ? {{28'd0}, _T_120} : _GEN_122;
  assign _GEN_125 = _T_40 ? 1'h0 : _GEN_113;
  assign _GEN_126 = _T_40 ? 1'h0 : _GEN_114;
  assign _GEN_127 = _T_40 ? 1'h0 : _GEN_115;
  assign _GEN_128 = _T_40 ? 1'h0 : _GEN_116;
  assign _GEN_129 = _T_40 ? 1'h0 : _GEN_117;
  assign _GEN_130 = _T_40 ? 1'h0 : _GEN_120;
  assign _GEN_133 = io_input_enable ? 1'h0 : 1'h1;
  assign _GEN_134 = io_input_enable ? _GEN_123 : 1'h0;
  assign _GEN_135 = io_input_enable ? _GEN_124 : 32'h1;
  assign _GEN_136 = io_input_enable ? _GEN_125 : 1'h0;
  assign _GEN_137 = io_input_enable ? _GEN_126 : 1'h0;
  assign _GEN_138 = io_input_enable ? _GEN_127 : 1'h0;
  assign _GEN_139 = io_input_enable ? _GEN_128 : 1'h0;
  assign _GEN_140 = io_input_enable ? _GEN_129 : 1'h0;
  assign _GEN_141 = io_input_enable ? _GEN_130 : 1'h0;
  assign _GEN_143 = io_input_enable ? _GEN_121 : 1'h0;
  assign _T_634 = ~ io_input_stageDone_0;
  assign _T_643 = io_input_stageDone_0 & _T_637;
  assign io_output_done = _T_91;
  assign io_output_stageEnable_0 = _GEN_136;
  assign io_output_stageEnable_1 = _GEN_137;
  assign io_output_stageEnable_2 = _GEN_138;
  assign io_output_stageEnable_3 = _GEN_139;
  assign io_output_stageEnable_4 = _GEN_140;
  assign io_output_rst_en = _T_102;
  assign io_output_ctr_inc = _T_643;
  assign deadState_io_input_set = _GEN_143;
  assign deadState_io_input_reset = _GEN_133;
  assign deadState_io_input_asyn_reset = _T_24;
  assign deadState_clock = clock;
  assign deadState_reset = reset;
  assign RetimeWrapper_io_flow = 1'h1;
  assign RetimeWrapper_io_in = reset;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_24 = RetimeWrapper_io_out;
  assign rstCtr_io_input_stop = 8'sh1;
  assign rstCtr_io_input_reset = _T_48;
  assign rstCtr_io_input_enable = _T_41;
  assign rstCtr_clock = clock;
  assign rstCtr_reset = reset;
  assign firstIterComplete_io_input_set = rstCtr_io_output_done;
  assign firstIterComplete_io_input_reset = _T_28;
  assign firstIterComplete_io_input_asyn_reset = _T_32;
  assign firstIterComplete_clock = clock;
  assign firstIterComplete_reset = reset;
  assign RetimeWrapper_1_io_flow = 1'h1;
  assign RetimeWrapper_1_io_in = reset;
  assign RetimeWrapper_1_clock = clock;
  assign RetimeWrapper_1_reset = reset;
  assign _T_28 = RetimeWrapper_1_io_out;
  assign RetimeWrapper_2_io_flow = 1'h1;
  assign RetimeWrapper_2_io_in = reset;
  assign RetimeWrapper_2_clock = clock;
  assign RetimeWrapper_2_reset = reset;
  assign _T_32 = RetimeWrapper_2_io_out;
  assign stateFF_io_input_0_data = _GEN_135;
  assign stateFF_io_input_0_init = 32'h1;
  assign stateFF_io_input_0_enable = 1'h1;
  assign stateFF_io_input_0_reset = _T_38;
  assign stateFF_clock = clock;
  assign stateFF_reset = reset;
  assign RetimeWrapper_3_io_flow = 1'h1;
  assign RetimeWrapper_3_io_in = io_input_rst;
  assign RetimeWrapper_3_clock = clock;
  assign RetimeWrapper_3_reset = reset;
  assign _T_38 = RetimeWrapper_3_io_out;
  assign RetimeWrapper_4_io_flow = 1'h1;
  assign RetimeWrapper_4_io_in = io_input_rst;
  assign RetimeWrapper_4_clock = clock;
  assign RetimeWrapper_4_reset = reset;
  assign _T_47 = RetimeWrapper_4_io_out;
  assign maxFF_io_input_0_data = io_input_numIter;
  assign maxFF_io_input_0_init = 32'h0;
  assign maxFF_io_input_0_enable = io_input_enable;
  assign maxFF_io_input_0_reset = _T_63;
  assign maxFF_clock = clock;
  assign maxFF_reset = reset;
  assign RetimeWrapper_5_io_flow = 1'h1;
  assign RetimeWrapper_5_io_in = io_input_rst;
  assign RetimeWrapper_5_clock = clock;
  assign RetimeWrapper_5_reset = reset;
  assign _T_63 = RetimeWrapper_5_io_out;
  assign RetimeWrapper_6_io_in = maxFF_io_output_data;
  assign RetimeWrapper_6_clock = clock;
  assign RetimeWrapper_6_reset = reset;
  assign max = RetimeWrapper_6_io_out;
  assign doneClear = _GEN_134;
  assign doneFF_0_io_input_set = io_input_stageDone_0;
  assign doneFF_0_io_input_reset = doneClear;
  assign doneFF_0_io_input_asyn_reset = _T_71;
  assign doneFF_0_clock = clock;
  assign doneFF_0_reset = reset;
  assign RetimeWrapper_7_io_flow = 1'h1;
  assign RetimeWrapper_7_io_in = io_input_rst;
  assign RetimeWrapper_7_clock = clock;
  assign RetimeWrapper_7_reset = reset;
  assign _T_71 = RetimeWrapper_7_io_out;
  assign doneFF_1_io_input_set = io_input_stageDone_1;
  assign doneFF_1_io_input_reset = doneClear;
  assign doneFF_1_io_input_asyn_reset = _T_75;
  assign doneFF_1_clock = clock;
  assign doneFF_1_reset = reset;
  assign RetimeWrapper_8_io_flow = 1'h1;
  assign RetimeWrapper_8_io_in = io_input_rst;
  assign RetimeWrapper_8_clock = clock;
  assign RetimeWrapper_8_reset = reset;
  assign _T_75 = RetimeWrapper_8_io_out;
  assign doneFF_2_io_input_set = io_input_stageDone_2;
  assign doneFF_2_io_input_reset = doneClear;
  assign doneFF_2_io_input_asyn_reset = _T_79;
  assign doneFF_2_clock = clock;
  assign doneFF_2_reset = reset;
  assign RetimeWrapper_9_io_flow = 1'h1;
  assign RetimeWrapper_9_io_in = io_input_rst;
  assign RetimeWrapper_9_clock = clock;
  assign RetimeWrapper_9_reset = reset;
  assign _T_79 = RetimeWrapper_9_io_out;
  assign doneFF_3_io_input_set = io_input_stageDone_3;
  assign doneFF_3_io_input_reset = doneClear;
  assign doneFF_3_io_input_asyn_reset = _T_83;
  assign doneFF_3_clock = clock;
  assign doneFF_3_reset = reset;
  assign RetimeWrapper_10_io_flow = 1'h1;
  assign RetimeWrapper_10_io_in = io_input_rst;
  assign RetimeWrapper_10_clock = clock;
  assign RetimeWrapper_10_reset = reset;
  assign _T_83 = RetimeWrapper_10_io_out;
  assign doneFF_4_io_input_set = io_input_stageDone_4;
  assign doneFF_4_io_input_reset = doneClear;
  assign doneFF_4_io_input_asyn_reset = _T_87;
  assign doneFF_4_clock = clock;
  assign doneFF_4_reset = reset;
  assign RetimeWrapper_11_io_flow = 1'h1;
  assign RetimeWrapper_11_io_in = io_input_rst;
  assign RetimeWrapper_11_clock = clock;
  assign RetimeWrapper_11_reset = reset;
  assign _T_87 = RetimeWrapper_11_io_out;
  assign ctr_io_input_stop = _T_89;
  assign ctr_io_input_stride = 32'sh0;
  assign ctr_io_input_reset = _T_96;
  assign ctr_io_input_enable = doneClear;
  assign ctr_io_input_saturate = 1'h1;
  assign ctr_clock = clock;
  assign ctr_reset = reset;
  assign RetimeWrapper_12_io_flow = 1'h1;
  assign RetimeWrapper_12_io_in = _T_92;
  assign RetimeWrapper_12_clock = clock;
  assign RetimeWrapper_12_reset = reset;
  assign _T_96 = RetimeWrapper_12_io_out;
  assign RetimeWrapper_13_io_flow = 1'h1;
  assign RetimeWrapper_13_io_in = _T_40;
  assign RetimeWrapper_13_clock = clock;
  assign RetimeWrapper_13_reset = reset;
  assign _T_102 = RetimeWrapper_13_io_out;
  assign cycsSinceDone_io_input_0_data = _GEN_32;
  assign cycsSinceDone_io_input_0_enable = _GEN_141;
  assign cycsSinceDone_io_input_0_reset = _T_91;
  assign cycsSinceDone_clock = clock;
  assign cycsSinceDone_reset = reset;
  assign RetimeWrapper_14_io_in = _T_484;
  assign RetimeWrapper_14_clock = clock;
  assign RetimeWrapper_14_reset = reset;
  assign _T_487 = _T_488;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_637 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_637 <= 1'h0;
    end else begin
      _T_637 <= _T_634;
    end
  end
endmodule
module RetimeWrapper_49(
  input        clock,
  input        reset,
  input  [3:0] io_in,
  output [3:0] io_out
);
  wire [3:0] sr_out;
  wire [3:0] sr_in;
  wire  sr_flow;
  wire  sr_reset;
  wire  sr_clock;
  RetimeShiftRegister #(.WIDTH(4), .STAGES(1)) sr (
    .out(sr_out),
    .in(sr_in),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out;
  assign sr_in = io_in;
  assign sr_flow = 1'h1;
  assign sr_reset = reset;
  assign sr_clock = clock;
endmodule
module NBufCtr(
  input        clock,
  input        reset,
  input        io_input_enable,
  output [3:0] io_output_count
);
  wire [3:0] _T_8;
  wire [4:0] _T_9;
  wire [3:0] _T_10;
  wire  _T_12;
  wire [4:0] _T_16;
  wire [4:0] _T_17;
  wire [3:0] _T_18;
  wire [3:0] _T_21;
  wire  _T_23;
  wire [4:0] _T_26;
  wire [4:0] _T_27;
  wire [3:0] _T_28;
  wire [3:0] _T_29;
  wire [3:0] _T_30;
  wire [3:0] _T_54;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire [3:0] RetimeWrapper_io_in;
  wire [3:0] RetimeWrapper_io_out;
  wire [3:0] _T_58;
  RetimeWrapper_49 RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_9 = _T_8 + 4'h0;
  assign _T_10 = _T_9[3:0];
  assign _T_12 = _T_10 >= 4'h5;
  assign _T_16 = _T_10 - 4'h5;
  assign _T_17 = $unsigned(_T_16);
  assign _T_18 = _T_17[3:0];
  assign _T_21 = _T_12 ? _T_18 : _T_10;
  assign _T_23 = _T_8 == 4'h0;
  assign _T_26 = _T_8 - 4'h1;
  assign _T_27 = $unsigned(_T_26);
  assign _T_28 = _T_27[3:0];
  assign _T_29 = _T_23 ? 4'h4 : _T_28;
  assign _T_30 = io_input_enable ? _T_29 : _T_8;
  assign _T_54 = reset ? 4'h0 : _T_30;
  assign io_output_count = _T_21;
  assign _T_8 = _T_58;
  assign RetimeWrapper_io_in = _T_54;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_58 = RetimeWrapper_io_out;
endmodule
module NBufCtr_1(
  input   clock,
  input   reset,
  input   io_input_enable
);
  wire [3:0] _T_8;
  wire  _T_25;
  wire [4:0] _T_28;
  wire [4:0] _T_29;
  wire [3:0] _T_30;
  wire [3:0] _T_31;
  wire [3:0] _T_32;
  wire [3:0] _T_55;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire [3:0] RetimeWrapper_io_in;
  wire [3:0] RetimeWrapper_io_out;
  wire [3:0] _T_59;
  RetimeWrapper_49 RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_25 = _T_8 == 4'h0;
  assign _T_28 = _T_8 - 4'h1;
  assign _T_29 = $unsigned(_T_28);
  assign _T_30 = _T_29[3:0];
  assign _T_31 = _T_25 ? 4'h4 : _T_30;
  assign _T_32 = io_input_enable ? _T_31 : _T_8;
  assign _T_55 = reset ? 4'h0 : _T_32;
  assign _T_8 = _T_59;
  assign RetimeWrapper_io_in = _T_55;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_59 = RetimeWrapper_io_out;
endmodule
module NBufCtr_2(
  input        clock,
  input        reset,
  input        io_input_enable,
  output [3:0] io_output_count
);
  wire [3:0] _T_8;
  wire [4:0] _T_10;
  wire [3:0] _T_11;
  wire  _T_13;
  wire [3:0] _T_14;
  wire [4:0] _T_16;
  wire [3:0] _T_17;
  wire [3:0] _T_18;
  wire [3:0] _T_19;
  wire [3:0] _T_23;
  wire  _T_25;
  wire [4:0] _T_28;
  wire [4:0] _T_29;
  wire [3:0] _T_30;
  wire [3:0] _T_31;
  wire [3:0] _T_32;
  wire [3:0] _T_55;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire [3:0] RetimeWrapper_io_in;
  wire [3:0] RetimeWrapper_io_out;
  wire [3:0] _T_59;
  RetimeWrapper_49 RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_10 = _T_8 + 4'h1;
  assign _T_11 = _T_10[3:0];
  assign _T_13 = _T_11 >= 4'h5;
  assign _T_14 = $signed(_T_8);
  assign _T_16 = $signed(_T_14) + $signed(-4'sh4);
  assign _T_17 = _T_16[3:0];
  assign _T_18 = $signed(_T_17);
  assign _T_19 = $unsigned(_T_18);
  assign _T_23 = _T_13 ? _T_19 : _T_11;
  assign _T_25 = _T_8 == 4'h0;
  assign _T_28 = _T_8 - 4'h1;
  assign _T_29 = $unsigned(_T_28);
  assign _T_30 = _T_29[3:0];
  assign _T_31 = _T_25 ? 4'h4 : _T_30;
  assign _T_32 = io_input_enable ? _T_31 : _T_8;
  assign _T_55 = reset ? 4'h0 : _T_32;
  assign io_output_count = _T_23;
  assign _T_8 = _T_59;
  assign RetimeWrapper_io_in = _T_55;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_59 = RetimeWrapper_io_out;
endmodule
module NBufCtr_3(
  input        clock,
  input        reset,
  input        io_input_enable,
  output [3:0] io_output_count
);
  wire [3:0] _T_8;
  wire [4:0] _T_10;
  wire [3:0] _T_11;
  wire  _T_13;
  wire [3:0] _T_14;
  wire [4:0] _T_16;
  wire [3:0] _T_17;
  wire [3:0] _T_18;
  wire [3:0] _T_19;
  wire [3:0] _T_23;
  wire  _T_25;
  wire [4:0] _T_28;
  wire [4:0] _T_29;
  wire [3:0] _T_30;
  wire [3:0] _T_31;
  wire [3:0] _T_32;
  wire [3:0] _T_55;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire [3:0] RetimeWrapper_io_in;
  wire [3:0] RetimeWrapper_io_out;
  wire [3:0] _T_59;
  RetimeWrapper_49 RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_10 = _T_8 + 4'h2;
  assign _T_11 = _T_10[3:0];
  assign _T_13 = _T_11 >= 4'h5;
  assign _T_14 = $signed(_T_8);
  assign _T_16 = $signed(_T_14) + $signed(-4'sh3);
  assign _T_17 = _T_16[3:0];
  assign _T_18 = $signed(_T_17);
  assign _T_19 = $unsigned(_T_18);
  assign _T_23 = _T_13 ? _T_19 : _T_11;
  assign _T_25 = _T_8 == 4'h0;
  assign _T_28 = _T_8 - 4'h1;
  assign _T_29 = $unsigned(_T_28);
  assign _T_30 = _T_29[3:0];
  assign _T_31 = _T_25 ? 4'h4 : _T_30;
  assign _T_32 = io_input_enable ? _T_31 : _T_8;
  assign _T_55 = reset ? 4'h0 : _T_32;
  assign io_output_count = _T_23;
  assign _T_8 = _T_59;
  assign RetimeWrapper_io_in = _T_55;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_59 = RetimeWrapper_io_out;
endmodule
module NBufCtr_4(
  input        clock,
  input        reset,
  input        io_input_enable,
  output [3:0] io_output_count
);
  wire [3:0] _T_8;
  wire [4:0] _T_10;
  wire [3:0] _T_11;
  wire  _T_13;
  wire [3:0] _T_14;
  wire [4:0] _T_16;
  wire [3:0] _T_17;
  wire [3:0] _T_18;
  wire [3:0] _T_19;
  wire [3:0] _T_23;
  wire  _T_25;
  wire [4:0] _T_28;
  wire [4:0] _T_29;
  wire [3:0] _T_30;
  wire [3:0] _T_31;
  wire [3:0] _T_32;
  wire [3:0] _T_55;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire [3:0] RetimeWrapper_io_in;
  wire [3:0] RetimeWrapper_io_out;
  wire [3:0] _T_59;
  RetimeWrapper_49 RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_10 = _T_8 + 4'h3;
  assign _T_11 = _T_10[3:0];
  assign _T_13 = _T_11 >= 4'h5;
  assign _T_14 = $signed(_T_8);
  assign _T_16 = $signed(_T_14) + $signed(-4'sh2);
  assign _T_17 = _T_16[3:0];
  assign _T_18 = $signed(_T_17);
  assign _T_19 = $unsigned(_T_18);
  assign _T_23 = _T_13 ? _T_19 : _T_11;
  assign _T_25 = _T_8 == 4'h0;
  assign _T_28 = _T_8 - 4'h1;
  assign _T_29 = $unsigned(_T_28);
  assign _T_30 = _T_29[3:0];
  assign _T_31 = _T_25 ? 4'h4 : _T_30;
  assign _T_32 = io_input_enable ? _T_31 : _T_8;
  assign _T_55 = reset ? 4'h0 : _T_32;
  assign io_output_count = _T_23;
  assign _T_8 = _T_59;
  assign RetimeWrapper_io_in = _T_55;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_59 = RetimeWrapper_io_out;
endmodule
module NBufCtr_5(
  input        clock,
  input        reset,
  input        io_input_enable,
  output [3:0] io_output_count
);
  wire [3:0] _T_8;
  wire [4:0] _T_10;
  wire [3:0] _T_11;
  wire  _T_13;
  wire [3:0] _T_14;
  wire [4:0] _T_16;
  wire [3:0] _T_17;
  wire [3:0] _T_18;
  wire [3:0] _T_19;
  wire [3:0] _T_23;
  wire  _T_25;
  wire [4:0] _T_28;
  wire [4:0] _T_29;
  wire [3:0] _T_30;
  wire [3:0] _T_31;
  wire [3:0] _T_32;
  wire [3:0] _T_55;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire [3:0] RetimeWrapper_io_in;
  wire [3:0] RetimeWrapper_io_out;
  wire [3:0] _T_59;
  RetimeWrapper_49 RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_10 = _T_8 + 4'h4;
  assign _T_11 = _T_10[3:0];
  assign _T_13 = _T_11 >= 4'h5;
  assign _T_14 = $signed(_T_8);
  assign _T_16 = $signed(_T_14) + $signed(-4'sh1);
  assign _T_17 = _T_16[3:0];
  assign _T_18 = $signed(_T_17);
  assign _T_19 = $unsigned(_T_18);
  assign _T_23 = _T_13 ? _T_19 : _T_11;
  assign _T_25 = _T_8 == 4'h0;
  assign _T_28 = _T_8 - 4'h1;
  assign _T_29 = $unsigned(_T_28);
  assign _T_30 = _T_29[3:0];
  assign _T_31 = _T_25 ? 4'h4 : _T_30;
  assign _T_32 = io_input_enable ? _T_31 : _T_8;
  assign _T_55 = reset ? 4'h0 : _T_32;
  assign io_output_count = _T_23;
  assign _T_8 = _T_59;
  assign RetimeWrapper_io_in = _T_55;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_59 = RetimeWrapper_io_out;
endmodule
module NBufFF(
  input         clock,
  input         reset,
  input         io_sEn_0,
  input         io_sEn_1,
  input         io_sEn_2,
  input         io_sEn_3,
  input         io_sEn_4,
  input         io_sDone_0,
  input         io_sDone_1,
  input         io_sDone_2,
  input         io_sDone_3,
  input         io_sDone_4,
  input  [31:0] io_input_0_data,
  input         io_input_0_enable,
  input         io_input_0_reset,
  output [31:0] io_output_1_data,
  output [31:0] io_output_2_data,
  output [31:0] io_output_4_data
);
  wire  ff_0_clock;
  wire  ff_0_reset;
  wire [31:0] ff_0_io_input_0_data;
  wire [31:0] ff_0_io_input_0_init;
  wire  ff_0_io_input_0_enable;
  wire  ff_0_io_input_0_reset;
  wire [31:0] ff_0_io_output_data;
  wire  ff_1_clock;
  wire  ff_1_reset;
  wire [31:0] ff_1_io_input_0_data;
  wire [31:0] ff_1_io_input_0_init;
  wire  ff_1_io_input_0_enable;
  wire  ff_1_io_input_0_reset;
  wire [31:0] ff_1_io_output_data;
  wire  ff_2_clock;
  wire  ff_2_reset;
  wire [31:0] ff_2_io_input_0_data;
  wire [31:0] ff_2_io_input_0_init;
  wire  ff_2_io_input_0_enable;
  wire  ff_2_io_input_0_reset;
  wire [31:0] ff_2_io_output_data;
  wire  ff_3_clock;
  wire  ff_3_reset;
  wire [31:0] ff_3_io_input_0_data;
  wire [31:0] ff_3_io_input_0_init;
  wire  ff_3_io_input_0_enable;
  wire  ff_3_io_input_0_reset;
  wire [31:0] ff_3_io_output_data;
  wire  ff_4_clock;
  wire  ff_4_reset;
  wire [31:0] ff_4_io_input_0_data;
  wire [31:0] ff_4_io_input_0_init;
  wire  ff_4_io_input_0_enable;
  wire  ff_4_io_input_0_reset;
  wire [31:0] ff_4_io_output_data;
  wire  sEn_latch_0_clock;
  wire  sEn_latch_0_reset;
  wire  sEn_latch_0_io_input_set;
  wire  sEn_latch_0_io_input_reset;
  wire  sEn_latch_0_io_input_asyn_reset;
  wire  sEn_latch_0_io_output_data;
  wire  sEn_latch_1_clock;
  wire  sEn_latch_1_reset;
  wire  sEn_latch_1_io_input_set;
  wire  sEn_latch_1_io_input_reset;
  wire  sEn_latch_1_io_input_asyn_reset;
  wire  sEn_latch_1_io_output_data;
  wire  sEn_latch_2_clock;
  wire  sEn_latch_2_reset;
  wire  sEn_latch_2_io_input_set;
  wire  sEn_latch_2_io_input_reset;
  wire  sEn_latch_2_io_input_asyn_reset;
  wire  sEn_latch_2_io_output_data;
  wire  sEn_latch_3_clock;
  wire  sEn_latch_3_reset;
  wire  sEn_latch_3_io_input_set;
  wire  sEn_latch_3_io_input_reset;
  wire  sEn_latch_3_io_input_asyn_reset;
  wire  sEn_latch_3_io_output_data;
  wire  sEn_latch_4_clock;
  wire  sEn_latch_4_reset;
  wire  sEn_latch_4_io_input_set;
  wire  sEn_latch_4_io_input_reset;
  wire  sEn_latch_4_io_input_asyn_reset;
  wire  sEn_latch_4_io_output_data;
  wire  sDone_latch_0_clock;
  wire  sDone_latch_0_reset;
  wire  sDone_latch_0_io_input_set;
  wire  sDone_latch_0_io_input_reset;
  wire  sDone_latch_0_io_input_asyn_reset;
  wire  sDone_latch_0_io_output_data;
  wire  sDone_latch_1_clock;
  wire  sDone_latch_1_reset;
  wire  sDone_latch_1_io_input_set;
  wire  sDone_latch_1_io_input_reset;
  wire  sDone_latch_1_io_input_asyn_reset;
  wire  sDone_latch_1_io_output_data;
  wire  sDone_latch_2_clock;
  wire  sDone_latch_2_reset;
  wire  sDone_latch_2_io_input_set;
  wire  sDone_latch_2_io_input_reset;
  wire  sDone_latch_2_io_input_asyn_reset;
  wire  sDone_latch_2_io_output_data;
  wire  sDone_latch_3_clock;
  wire  sDone_latch_3_reset;
  wire  sDone_latch_3_io_input_set;
  wire  sDone_latch_3_io_input_reset;
  wire  sDone_latch_3_io_input_asyn_reset;
  wire  sDone_latch_3_io_output_data;
  wire  sDone_latch_4_clock;
  wire  sDone_latch_4_reset;
  wire  sDone_latch_4_io_input_set;
  wire  sDone_latch_4_io_input_reset;
  wire  sDone_latch_4_io_input_asyn_reset;
  wire  sDone_latch_4_io_output_data;
  wire  swap;
  wire  _T_20;
  wire  _T_21;
  wire  _T_22;
  wire  _T_23;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire  RetimeWrapper_io_flow;
  wire  RetimeWrapper_io_in;
  wire  RetimeWrapper_io_out;
  wire  _T_27;
  wire  _T_28;
  wire  _T_29;
  wire  RetimeWrapper_1_clock;
  wire  RetimeWrapper_1_reset;
  wire  RetimeWrapper_1_io_flow;
  wire  RetimeWrapper_1_io_in;
  wire  RetimeWrapper_1_io_out;
  wire  _T_33;
  wire  _T_34;
  wire  RetimeWrapper_2_clock;
  wire  RetimeWrapper_2_reset;
  wire  RetimeWrapper_2_io_flow;
  wire  RetimeWrapper_2_io_in;
  wire  RetimeWrapper_2_io_out;
  wire  _T_38;
  wire  RetimeWrapper_3_clock;
  wire  RetimeWrapper_3_reset;
  wire  RetimeWrapper_3_io_flow;
  wire  RetimeWrapper_3_io_in;
  wire  RetimeWrapper_3_io_out;
  wire  _T_42;
  wire  _T_43;
  wire  RetimeWrapper_4_clock;
  wire  RetimeWrapper_4_reset;
  wire  RetimeWrapper_4_io_flow;
  wire  RetimeWrapper_4_io_in;
  wire  RetimeWrapper_4_io_out;
  wire  _T_47;
  wire  _T_48;
  wire  _T_49;
  wire  _T_50;
  wire  _T_51;
  wire  RetimeWrapper_5_clock;
  wire  RetimeWrapper_5_reset;
  wire  RetimeWrapper_5_io_flow;
  wire  RetimeWrapper_5_io_in;
  wire  RetimeWrapper_5_io_out;
  wire  _T_55;
  wire  _T_56;
  wire  _T_57;
  wire  RetimeWrapper_6_clock;
  wire  RetimeWrapper_6_reset;
  wire  RetimeWrapper_6_io_flow;
  wire  RetimeWrapper_6_io_in;
  wire  RetimeWrapper_6_io_out;
  wire  _T_61;
  wire  _T_62;
  wire  RetimeWrapper_7_clock;
  wire  RetimeWrapper_7_reset;
  wire  RetimeWrapper_7_io_flow;
  wire  RetimeWrapper_7_io_in;
  wire  RetimeWrapper_7_io_out;
  wire  _T_66;
  wire  RetimeWrapper_8_clock;
  wire  RetimeWrapper_8_reset;
  wire  RetimeWrapper_8_io_flow;
  wire  RetimeWrapper_8_io_in;
  wire  RetimeWrapper_8_io_out;
  wire  _T_70;
  wire  _T_71;
  wire  RetimeWrapper_9_clock;
  wire  RetimeWrapper_9_reset;
  wire  RetimeWrapper_9_io_flow;
  wire  RetimeWrapper_9_io_in;
  wire  RetimeWrapper_9_io_out;
  wire  _T_75;
  wire  _T_76;
  wire  _T_77;
  wire  _T_78;
  wire  _T_79;
  wire  RetimeWrapper_10_clock;
  wire  RetimeWrapper_10_reset;
  wire  RetimeWrapper_10_io_flow;
  wire  RetimeWrapper_10_io_in;
  wire  RetimeWrapper_10_io_out;
  wire  _T_83;
  wire  _T_84;
  wire  _T_85;
  wire  RetimeWrapper_11_clock;
  wire  RetimeWrapper_11_reset;
  wire  RetimeWrapper_11_io_flow;
  wire  RetimeWrapper_11_io_in;
  wire  RetimeWrapper_11_io_out;
  wire  _T_89;
  wire  _T_90;
  wire  RetimeWrapper_12_clock;
  wire  RetimeWrapper_12_reset;
  wire  RetimeWrapper_12_io_flow;
  wire  RetimeWrapper_12_io_in;
  wire  RetimeWrapper_12_io_out;
  wire  _T_94;
  wire  RetimeWrapper_13_clock;
  wire  RetimeWrapper_13_reset;
  wire  RetimeWrapper_13_io_flow;
  wire  RetimeWrapper_13_io_in;
  wire  RetimeWrapper_13_io_out;
  wire  _T_98;
  wire  _T_99;
  wire  RetimeWrapper_14_clock;
  wire  RetimeWrapper_14_reset;
  wire  RetimeWrapper_14_io_flow;
  wire  RetimeWrapper_14_io_in;
  wire  RetimeWrapper_14_io_out;
  wire  _T_103;
  wire  _T_104;
  wire  _T_105;
  wire  _T_106;
  wire  _T_107;
  wire  RetimeWrapper_15_clock;
  wire  RetimeWrapper_15_reset;
  wire  RetimeWrapper_15_io_flow;
  wire  RetimeWrapper_15_io_in;
  wire  RetimeWrapper_15_io_out;
  wire  _T_111;
  wire  _T_112;
  wire  _T_113;
  wire  RetimeWrapper_16_clock;
  wire  RetimeWrapper_16_reset;
  wire  RetimeWrapper_16_io_flow;
  wire  RetimeWrapper_16_io_in;
  wire  RetimeWrapper_16_io_out;
  wire  _T_117;
  wire  _T_118;
  wire  RetimeWrapper_17_clock;
  wire  RetimeWrapper_17_reset;
  wire  RetimeWrapper_17_io_flow;
  wire  RetimeWrapper_17_io_in;
  wire  RetimeWrapper_17_io_out;
  wire  _T_122;
  wire  RetimeWrapper_18_clock;
  wire  RetimeWrapper_18_reset;
  wire  RetimeWrapper_18_io_flow;
  wire  RetimeWrapper_18_io_in;
  wire  RetimeWrapper_18_io_out;
  wire  _T_126;
  wire  _T_127;
  wire  RetimeWrapper_19_clock;
  wire  RetimeWrapper_19_reset;
  wire  RetimeWrapper_19_io_flow;
  wire  RetimeWrapper_19_io_in;
  wire  RetimeWrapper_19_io_out;
  wire  _T_131;
  wire  _T_132;
  wire  _T_133;
  wire  _T_134;
  wire  _T_135;
  wire  RetimeWrapper_20_clock;
  wire  RetimeWrapper_20_reset;
  wire  RetimeWrapper_20_io_flow;
  wire  RetimeWrapper_20_io_in;
  wire  RetimeWrapper_20_io_out;
  wire  _T_139;
  wire  _T_140;
  wire  _T_141;
  wire  RetimeWrapper_21_clock;
  wire  RetimeWrapper_21_reset;
  wire  RetimeWrapper_21_io_flow;
  wire  RetimeWrapper_21_io_in;
  wire  RetimeWrapper_21_io_out;
  wire  _T_145;
  wire  _T_146;
  wire  RetimeWrapper_22_clock;
  wire  RetimeWrapper_22_reset;
  wire  RetimeWrapper_22_io_flow;
  wire  RetimeWrapper_22_io_in;
  wire  RetimeWrapper_22_io_out;
  wire  _T_150;
  wire  RetimeWrapper_23_clock;
  wire  RetimeWrapper_23_reset;
  wire  RetimeWrapper_23_io_flow;
  wire  RetimeWrapper_23_io_in;
  wire  RetimeWrapper_23_io_out;
  wire  _T_154;
  wire  _T_155;
  wire  RetimeWrapper_24_clock;
  wire  RetimeWrapper_24_reset;
  wire  RetimeWrapper_24_io_flow;
  wire  RetimeWrapper_24_io_in;
  wire  RetimeWrapper_24_io_out;
  wire  _T_159;
  wire  _T_160;
  wire  _T_161;
  wire  _T_162;
  wire  anyEnabled;
  wire  _T_163;
  wire  _T_164;
  wire  _T_165;
  wire  _T_166;
  wire  _T_167;
  wire  _T_168;
  wire  _T_169;
  wire  _T_170;
  wire  _T_171;
  wire  _T_172;
  wire  _T_173;
  wire  _T_174;
  wire  _T_175;
  wire  _T_176;
  wire  _T_177;
  wire  _T_178;
  reg  _T_181;
  reg [31:0] _RAND_0;
  wire  _T_187;
  wire  statesIn_0_clock;
  wire  statesIn_0_reset;
  wire  statesIn_0_io_input_enable;
  wire [3:0] statesIn_0_io_output_count;
  wire  statesOut_0_clock;
  wire  statesOut_0_reset;
  wire  statesOut_0_io_input_enable;
  wire  statesOut_1_clock;
  wire  statesOut_1_reset;
  wire  statesOut_1_io_input_enable;
  wire [3:0] statesOut_1_io_output_count;
  wire  statesOut_2_clock;
  wire  statesOut_2_reset;
  wire  statesOut_2_io_input_enable;
  wire [3:0] statesOut_2_io_output_count;
  wire  statesOut_3_clock;
  wire  statesOut_3_reset;
  wire  statesOut_3_io_input_enable;
  wire [3:0] statesOut_3_io_output_count;
  wire  statesOut_4_clock;
  wire  statesOut_4_reset;
  wire  statesOut_4_io_input_enable;
  wire [3:0] statesOut_4_io_output_count;
  wire  _T_195;
  wire [31:0] _T_197_data;
  wire  _T_197_enable;
  wire  _T_197_reset;
  wire  _T_198;
  wire  _T_201;
  wire [31:0] _T_203_data;
  wire  _T_203_enable;
  wire  _T_203_reset;
  wire  _T_204;
  wire  _T_207;
  wire [31:0] _T_209_data;
  wire  _T_209_enable;
  wire  _T_209_reset;
  wire  _T_210;
  wire  _T_213;
  wire [31:0] _T_215_data;
  wire  _T_215_enable;
  wire  _T_215_reset;
  wire  _T_216;
  wire  _T_219;
  wire [31:0] _T_221_data;
  wire  _T_221_enable;
  wire  _T_221_reset;
  wire  _T_222;
  wire  _T_262;
  wire  _T_264;
  wire  _T_266;
  wire  _T_268;
  wire  _T_270;
  wire [31:0] _T_273_0;
  wire [31:0] _T_273_1;
  wire [31:0] _T_273_2;
  wire [31:0] _T_273_3;
  wire [31:0] _T_273_4;
  wire [31:0] _T_283;
  wire [31:0] _T_285;
  wire [31:0] _T_287;
  wire [31:0] _T_289;
  wire [31:0] _T_291;
  wire [31:0] _T_292;
  wire [31:0] _T_293;
  wire [31:0] _T_294;
  wire [31:0] _T_295;
  wire [31:0] _T_297;
  wire  _T_299;
  wire  _T_301;
  wire  _T_303;
  wire  _T_305;
  wire  _T_307;
  wire [31:0] _T_310_0;
  wire [31:0] _T_310_1;
  wire [31:0] _T_310_2;
  wire [31:0] _T_310_3;
  wire [31:0] _T_310_4;
  wire [31:0] _T_320;
  wire [31:0] _T_322;
  wire [31:0] _T_324;
  wire [31:0] _T_326;
  wire [31:0] _T_328;
  wire [31:0] _T_329;
  wire [31:0] _T_330;
  wire [31:0] _T_331;
  wire [31:0] _T_332;
  wire [31:0] _T_334;
  wire  _T_373;
  wire  _T_375;
  wire  _T_377;
  wire  _T_379;
  wire  _T_381;
  wire [31:0] _T_384_0;
  wire [31:0] _T_384_1;
  wire [31:0] _T_384_2;
  wire [31:0] _T_384_3;
  wire [31:0] _T_384_4;
  wire [31:0] _T_394;
  wire [31:0] _T_396;
  wire [31:0] _T_398;
  wire [31:0] _T_400;
  wire [31:0] _T_402;
  wire [31:0] _T_403;
  wire [31:0] _T_404;
  wire [31:0] _T_405;
  wire [31:0] _T_406;
  wire [31:0] _T_408;
  FF_1 ff_0 (
    .clock(ff_0_clock),
    .reset(ff_0_reset),
    .io_input_0_data(ff_0_io_input_0_data),
    .io_input_0_init(ff_0_io_input_0_init),
    .io_input_0_enable(ff_0_io_input_0_enable),
    .io_input_0_reset(ff_0_io_input_0_reset),
    .io_output_data(ff_0_io_output_data)
  );
  FF_1 ff_1 (
    .clock(ff_1_clock),
    .reset(ff_1_reset),
    .io_input_0_data(ff_1_io_input_0_data),
    .io_input_0_init(ff_1_io_input_0_init),
    .io_input_0_enable(ff_1_io_input_0_enable),
    .io_input_0_reset(ff_1_io_input_0_reset),
    .io_output_data(ff_1_io_output_data)
  );
  FF_1 ff_2 (
    .clock(ff_2_clock),
    .reset(ff_2_reset),
    .io_input_0_data(ff_2_io_input_0_data),
    .io_input_0_init(ff_2_io_input_0_init),
    .io_input_0_enable(ff_2_io_input_0_enable),
    .io_input_0_reset(ff_2_io_input_0_reset),
    .io_output_data(ff_2_io_output_data)
  );
  FF_1 ff_3 (
    .clock(ff_3_clock),
    .reset(ff_3_reset),
    .io_input_0_data(ff_3_io_input_0_data),
    .io_input_0_init(ff_3_io_input_0_init),
    .io_input_0_enable(ff_3_io_input_0_enable),
    .io_input_0_reset(ff_3_io_input_0_reset),
    .io_output_data(ff_3_io_output_data)
  );
  FF_1 ff_4 (
    .clock(ff_4_clock),
    .reset(ff_4_reset),
    .io_input_0_data(ff_4_io_input_0_data),
    .io_input_0_init(ff_4_io_input_0_init),
    .io_input_0_enable(ff_4_io_input_0_enable),
    .io_input_0_reset(ff_4_io_input_0_reset),
    .io_output_data(ff_4_io_output_data)
  );
  SRFF sEn_latch_0 (
    .clock(sEn_latch_0_clock),
    .reset(sEn_latch_0_reset),
    .io_input_set(sEn_latch_0_io_input_set),
    .io_input_reset(sEn_latch_0_io_input_reset),
    .io_input_asyn_reset(sEn_latch_0_io_input_asyn_reset),
    .io_output_data(sEn_latch_0_io_output_data)
  );
  SRFF sEn_latch_1 (
    .clock(sEn_latch_1_clock),
    .reset(sEn_latch_1_reset),
    .io_input_set(sEn_latch_1_io_input_set),
    .io_input_reset(sEn_latch_1_io_input_reset),
    .io_input_asyn_reset(sEn_latch_1_io_input_asyn_reset),
    .io_output_data(sEn_latch_1_io_output_data)
  );
  SRFF sEn_latch_2 (
    .clock(sEn_latch_2_clock),
    .reset(sEn_latch_2_reset),
    .io_input_set(sEn_latch_2_io_input_set),
    .io_input_reset(sEn_latch_2_io_input_reset),
    .io_input_asyn_reset(sEn_latch_2_io_input_asyn_reset),
    .io_output_data(sEn_latch_2_io_output_data)
  );
  SRFF sEn_latch_3 (
    .clock(sEn_latch_3_clock),
    .reset(sEn_latch_3_reset),
    .io_input_set(sEn_latch_3_io_input_set),
    .io_input_reset(sEn_latch_3_io_input_reset),
    .io_input_asyn_reset(sEn_latch_3_io_input_asyn_reset),
    .io_output_data(sEn_latch_3_io_output_data)
  );
  SRFF sEn_latch_4 (
    .clock(sEn_latch_4_clock),
    .reset(sEn_latch_4_reset),
    .io_input_set(sEn_latch_4_io_input_set),
    .io_input_reset(sEn_latch_4_io_input_reset),
    .io_input_asyn_reset(sEn_latch_4_io_input_asyn_reset),
    .io_output_data(sEn_latch_4_io_output_data)
  );
  SRFF sDone_latch_0 (
    .clock(sDone_latch_0_clock),
    .reset(sDone_latch_0_reset),
    .io_input_set(sDone_latch_0_io_input_set),
    .io_input_reset(sDone_latch_0_io_input_reset),
    .io_input_asyn_reset(sDone_latch_0_io_input_asyn_reset),
    .io_output_data(sDone_latch_0_io_output_data)
  );
  SRFF sDone_latch_1 (
    .clock(sDone_latch_1_clock),
    .reset(sDone_latch_1_reset),
    .io_input_set(sDone_latch_1_io_input_set),
    .io_input_reset(sDone_latch_1_io_input_reset),
    .io_input_asyn_reset(sDone_latch_1_io_input_asyn_reset),
    .io_output_data(sDone_latch_1_io_output_data)
  );
  SRFF sDone_latch_2 (
    .clock(sDone_latch_2_clock),
    .reset(sDone_latch_2_reset),
    .io_input_set(sDone_latch_2_io_input_set),
    .io_input_reset(sDone_latch_2_io_input_reset),
    .io_input_asyn_reset(sDone_latch_2_io_input_asyn_reset),
    .io_output_data(sDone_latch_2_io_output_data)
  );
  SRFF sDone_latch_3 (
    .clock(sDone_latch_3_clock),
    .reset(sDone_latch_3_reset),
    .io_input_set(sDone_latch_3_io_input_set),
    .io_input_reset(sDone_latch_3_io_input_reset),
    .io_input_asyn_reset(sDone_latch_3_io_input_asyn_reset),
    .io_output_data(sDone_latch_3_io_output_data)
  );
  SRFF sDone_latch_4 (
    .clock(sDone_latch_4_clock),
    .reset(sDone_latch_4_reset),
    .io_input_set(sDone_latch_4_io_input_set),
    .io_input_reset(sDone_latch_4_io_input_reset),
    .io_input_asyn_reset(sDone_latch_4_io_input_asyn_reset),
    .io_output_data(sDone_latch_4_io_output_data)
  );
  RetimeWrapper RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 (
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 (
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 (
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 (
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 (
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 (
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 (
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper RetimeWrapper_8 (
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper RetimeWrapper_9 (
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper RetimeWrapper_10 (
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper RetimeWrapper_11 (
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper RetimeWrapper_12 (
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper RetimeWrapper_13 (
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper RetimeWrapper_14 (
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper RetimeWrapper_15 (
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper RetimeWrapper_16 (
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper RetimeWrapper_17 (
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper RetimeWrapper_18 (
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper RetimeWrapper_19 (
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper RetimeWrapper_20 (
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper RetimeWrapper_21 (
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper RetimeWrapper_22 (
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper RetimeWrapper_23 (
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper RetimeWrapper_24 (
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  NBufCtr statesIn_0 (
    .clock(statesIn_0_clock),
    .reset(statesIn_0_reset),
    .io_input_enable(statesIn_0_io_input_enable),
    .io_output_count(statesIn_0_io_output_count)
  );
  NBufCtr_1 statesOut_0 (
    .clock(statesOut_0_clock),
    .reset(statesOut_0_reset),
    .io_input_enable(statesOut_0_io_input_enable)
  );
  NBufCtr_2 statesOut_1 (
    .clock(statesOut_1_clock),
    .reset(statesOut_1_reset),
    .io_input_enable(statesOut_1_io_input_enable),
    .io_output_count(statesOut_1_io_output_count)
  );
  NBufCtr_3 statesOut_2 (
    .clock(statesOut_2_clock),
    .reset(statesOut_2_reset),
    .io_input_enable(statesOut_2_io_input_enable),
    .io_output_count(statesOut_2_io_output_count)
  );
  NBufCtr_4 statesOut_3 (
    .clock(statesOut_3_clock),
    .reset(statesOut_3_reset),
    .io_input_enable(statesOut_3_io_input_enable),
    .io_output_count(statesOut_3_io_output_count)
  );
  NBufCtr_5 statesOut_4 (
    .clock(statesOut_4_clock),
    .reset(statesOut_4_reset),
    .io_input_enable(statesOut_4_io_input_enable),
    .io_output_count(statesOut_4_io_output_count)
  );
  assign _T_20 = ~ io_sDone_0;
  assign _T_21 = io_sEn_0 & _T_20;
  assign _T_22 = io_sEn_0 & io_sDone_0;
  assign _T_23 = ~ io_sEn_0;
  assign _T_28 = _T_22 & _T_27;
  assign _T_29 = _T_21 | _T_28;
  assign _T_34 = swap | _T_33;
  assign _T_43 = swap | _T_42;
  assign _T_48 = ~ io_sDone_1;
  assign _T_49 = io_sEn_1 & _T_48;
  assign _T_50 = io_sEn_1 & io_sDone_1;
  assign _T_51 = ~ io_sEn_1;
  assign _T_56 = _T_50 & _T_55;
  assign _T_57 = _T_49 | _T_56;
  assign _T_62 = swap | _T_61;
  assign _T_71 = swap | _T_70;
  assign _T_76 = ~ io_sDone_2;
  assign _T_77 = io_sEn_2 & _T_76;
  assign _T_78 = io_sEn_2 & io_sDone_2;
  assign _T_79 = ~ io_sEn_2;
  assign _T_84 = _T_78 & _T_83;
  assign _T_85 = _T_77 | _T_84;
  assign _T_90 = swap | _T_89;
  assign _T_99 = swap | _T_98;
  assign _T_104 = ~ io_sDone_3;
  assign _T_105 = io_sEn_3 & _T_104;
  assign _T_106 = io_sEn_3 & io_sDone_3;
  assign _T_107 = ~ io_sEn_3;
  assign _T_112 = _T_106 & _T_111;
  assign _T_113 = _T_105 | _T_112;
  assign _T_118 = swap | _T_117;
  assign _T_127 = swap | _T_126;
  assign _T_132 = ~ io_sDone_4;
  assign _T_133 = io_sEn_4 & _T_132;
  assign _T_134 = io_sEn_4 & io_sDone_4;
  assign _T_135 = ~ io_sEn_4;
  assign _T_140 = _T_134 & _T_139;
  assign _T_141 = _T_133 | _T_140;
  assign _T_146 = swap | _T_145;
  assign _T_155 = swap | _T_154;
  assign _T_160 = sEn_latch_0_io_output_data | sEn_latch_1_io_output_data;
  assign _T_161 = _T_160 | sEn_latch_2_io_output_data;
  assign _T_162 = _T_161 | sEn_latch_3_io_output_data;
  assign anyEnabled = _T_162 | sEn_latch_4_io_output_data;
  assign _T_163 = sDone_latch_0_io_output_data | io_sDone_0;
  assign _T_164 = sEn_latch_0_io_output_data == _T_163;
  assign _T_165 = sDone_latch_1_io_output_data | io_sDone_1;
  assign _T_166 = sEn_latch_1_io_output_data == _T_165;
  assign _T_167 = sDone_latch_2_io_output_data | io_sDone_2;
  assign _T_168 = sEn_latch_2_io_output_data == _T_167;
  assign _T_169 = sDone_latch_3_io_output_data | io_sDone_3;
  assign _T_170 = sEn_latch_3_io_output_data == _T_169;
  assign _T_171 = sDone_latch_4_io_output_data | io_sDone_4;
  assign _T_172 = sEn_latch_4_io_output_data == _T_171;
  assign _T_173 = _T_164 & _T_166;
  assign _T_174 = _T_173 & _T_168;
  assign _T_175 = _T_174 & _T_170;
  assign _T_176 = _T_175 & _T_172;
  assign _T_177 = _T_176 & anyEnabled;
  assign _T_178 = ~ _T_177;
  assign _T_187 = _T_177 & _T_181;
  assign _T_195 = statesIn_0_io_output_count == 4'h0;
  assign _T_198 = io_input_0_enable & _T_195;
  assign _T_201 = statesIn_0_io_output_count == 4'h1;
  assign _T_204 = io_input_0_enable & _T_201;
  assign _T_207 = statesIn_0_io_output_count == 4'h2;
  assign _T_210 = io_input_0_enable & _T_207;
  assign _T_213 = statesIn_0_io_output_count == 4'h3;
  assign _T_216 = io_input_0_enable & _T_213;
  assign _T_219 = statesIn_0_io_output_count == 4'h4;
  assign _T_222 = io_input_0_enable & _T_219;
  assign _T_262 = statesOut_1_io_output_count == 4'h0;
  assign _T_264 = statesOut_1_io_output_count == 4'h1;
  assign _T_266 = statesOut_1_io_output_count == 4'h2;
  assign _T_268 = statesOut_1_io_output_count == 4'h3;
  assign _T_270 = statesOut_1_io_output_count == 4'h4;
  assign _T_283 = _T_262 ? _T_273_0 : 32'h0;
  assign _T_285 = _T_264 ? _T_273_1 : 32'h0;
  assign _T_287 = _T_266 ? _T_273_2 : 32'h0;
  assign _T_289 = _T_268 ? _T_273_3 : 32'h0;
  assign _T_291 = _T_270 ? _T_273_4 : 32'h0;
  assign _T_292 = _T_283 | _T_285;
  assign _T_293 = _T_292 | _T_287;
  assign _T_294 = _T_293 | _T_289;
  assign _T_295 = _T_294 | _T_291;
  assign _T_299 = statesOut_2_io_output_count == 4'h0;
  assign _T_301 = statesOut_2_io_output_count == 4'h1;
  assign _T_303 = statesOut_2_io_output_count == 4'h2;
  assign _T_305 = statesOut_2_io_output_count == 4'h3;
  assign _T_307 = statesOut_2_io_output_count == 4'h4;
  assign _T_320 = _T_299 ? _T_310_0 : 32'h0;
  assign _T_322 = _T_301 ? _T_310_1 : 32'h0;
  assign _T_324 = _T_303 ? _T_310_2 : 32'h0;
  assign _T_326 = _T_305 ? _T_310_3 : 32'h0;
  assign _T_328 = _T_307 ? _T_310_4 : 32'h0;
  assign _T_329 = _T_320 | _T_322;
  assign _T_330 = _T_329 | _T_324;
  assign _T_331 = _T_330 | _T_326;
  assign _T_332 = _T_331 | _T_328;
  assign _T_373 = statesOut_4_io_output_count == 4'h0;
  assign _T_375 = statesOut_4_io_output_count == 4'h1;
  assign _T_377 = statesOut_4_io_output_count == 4'h2;
  assign _T_379 = statesOut_4_io_output_count == 4'h3;
  assign _T_381 = statesOut_4_io_output_count == 4'h4;
  assign _T_394 = _T_373 ? _T_384_0 : 32'h0;
  assign _T_396 = _T_375 ? _T_384_1 : 32'h0;
  assign _T_398 = _T_377 ? _T_384_2 : 32'h0;
  assign _T_400 = _T_379 ? _T_384_3 : 32'h0;
  assign _T_402 = _T_381 ? _T_384_4 : 32'h0;
  assign _T_403 = _T_394 | _T_396;
  assign _T_404 = _T_403 | _T_398;
  assign _T_405 = _T_404 | _T_400;
  assign _T_406 = _T_405 | _T_402;
  assign io_output_1_data = _T_297;
  assign io_output_2_data = _T_334;
  assign io_output_4_data = _T_408;
  assign ff_0_io_input_0_data = _T_197_data;
  assign ff_0_io_input_0_init = 32'h0;
  assign ff_0_io_input_0_enable = _T_197_enable;
  assign ff_0_io_input_0_reset = _T_197_reset;
  assign ff_0_clock = clock;
  assign ff_0_reset = reset;
  assign ff_1_io_input_0_data = _T_203_data;
  assign ff_1_io_input_0_init = 32'h0;
  assign ff_1_io_input_0_enable = _T_203_enable;
  assign ff_1_io_input_0_reset = _T_203_reset;
  assign ff_1_clock = clock;
  assign ff_1_reset = reset;
  assign ff_2_io_input_0_data = _T_209_data;
  assign ff_2_io_input_0_init = 32'h0;
  assign ff_2_io_input_0_enable = _T_209_enable;
  assign ff_2_io_input_0_reset = _T_209_reset;
  assign ff_2_clock = clock;
  assign ff_2_reset = reset;
  assign ff_3_io_input_0_data = _T_215_data;
  assign ff_3_io_input_0_init = 32'h0;
  assign ff_3_io_input_0_enable = _T_215_enable;
  assign ff_3_io_input_0_reset = _T_215_reset;
  assign ff_3_clock = clock;
  assign ff_3_reset = reset;
  assign ff_4_io_input_0_data = _T_221_data;
  assign ff_4_io_input_0_init = 32'h0;
  assign ff_4_io_input_0_enable = _T_221_enable;
  assign ff_4_io_input_0_reset = _T_221_reset;
  assign ff_4_clock = clock;
  assign ff_4_reset = reset;
  assign sEn_latch_0_io_input_set = _T_29;
  assign sEn_latch_0_io_input_reset = _T_34;
  assign sEn_latch_0_io_input_asyn_reset = _T_38;
  assign sEn_latch_0_clock = clock;
  assign sEn_latch_0_reset = reset;
  assign sEn_latch_1_io_input_set = _T_57;
  assign sEn_latch_1_io_input_reset = _T_62;
  assign sEn_latch_1_io_input_asyn_reset = _T_66;
  assign sEn_latch_1_clock = clock;
  assign sEn_latch_1_reset = reset;
  assign sEn_latch_2_io_input_set = _T_85;
  assign sEn_latch_2_io_input_reset = _T_90;
  assign sEn_latch_2_io_input_asyn_reset = _T_94;
  assign sEn_latch_2_clock = clock;
  assign sEn_latch_2_reset = reset;
  assign sEn_latch_3_io_input_set = _T_113;
  assign sEn_latch_3_io_input_reset = _T_118;
  assign sEn_latch_3_io_input_asyn_reset = _T_122;
  assign sEn_latch_3_clock = clock;
  assign sEn_latch_3_reset = reset;
  assign sEn_latch_4_io_input_set = _T_141;
  assign sEn_latch_4_io_input_reset = _T_146;
  assign sEn_latch_4_io_input_asyn_reset = _T_150;
  assign sEn_latch_4_clock = clock;
  assign sEn_latch_4_reset = reset;
  assign sDone_latch_0_io_input_set = io_sDone_0;
  assign sDone_latch_0_io_input_reset = _T_43;
  assign sDone_latch_0_io_input_asyn_reset = _T_47;
  assign sDone_latch_0_clock = clock;
  assign sDone_latch_0_reset = reset;
  assign sDone_latch_1_io_input_set = io_sDone_1;
  assign sDone_latch_1_io_input_reset = _T_71;
  assign sDone_latch_1_io_input_asyn_reset = _T_75;
  assign sDone_latch_1_clock = clock;
  assign sDone_latch_1_reset = reset;
  assign sDone_latch_2_io_input_set = io_sDone_2;
  assign sDone_latch_2_io_input_reset = _T_99;
  assign sDone_latch_2_io_input_asyn_reset = _T_103;
  assign sDone_latch_2_clock = clock;
  assign sDone_latch_2_reset = reset;
  assign sDone_latch_3_io_input_set = io_sDone_3;
  assign sDone_latch_3_io_input_reset = _T_127;
  assign sDone_latch_3_io_input_asyn_reset = _T_131;
  assign sDone_latch_3_clock = clock;
  assign sDone_latch_3_reset = reset;
  assign sDone_latch_4_io_input_set = io_sDone_4;
  assign sDone_latch_4_io_input_reset = _T_155;
  assign sDone_latch_4_io_input_asyn_reset = _T_159;
  assign sDone_latch_4_clock = clock;
  assign sDone_latch_4_reset = reset;
  assign swap = _T_187;
  assign RetimeWrapper_io_flow = 1'h1;
  assign RetimeWrapper_io_in = _T_23;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_27 = RetimeWrapper_io_out;
  assign RetimeWrapper_1_io_flow = 1'h1;
  assign RetimeWrapper_1_io_in = swap;
  assign RetimeWrapper_1_clock = clock;
  assign RetimeWrapper_1_reset = reset;
  assign _T_33 = RetimeWrapper_1_io_out;
  assign RetimeWrapper_2_io_flow = 1'h1;
  assign RetimeWrapper_2_io_in = reset;
  assign RetimeWrapper_2_clock = clock;
  assign RetimeWrapper_2_reset = reset;
  assign _T_38 = RetimeWrapper_2_io_out;
  assign RetimeWrapper_3_io_flow = 1'h1;
  assign RetimeWrapper_3_io_in = swap;
  assign RetimeWrapper_3_clock = clock;
  assign RetimeWrapper_3_reset = reset;
  assign _T_42 = RetimeWrapper_3_io_out;
  assign RetimeWrapper_4_io_flow = 1'h1;
  assign RetimeWrapper_4_io_in = reset;
  assign RetimeWrapper_4_clock = clock;
  assign RetimeWrapper_4_reset = reset;
  assign _T_47 = RetimeWrapper_4_io_out;
  assign RetimeWrapper_5_io_flow = 1'h1;
  assign RetimeWrapper_5_io_in = _T_51;
  assign RetimeWrapper_5_clock = clock;
  assign RetimeWrapper_5_reset = reset;
  assign _T_55 = RetimeWrapper_5_io_out;
  assign RetimeWrapper_6_io_flow = 1'h1;
  assign RetimeWrapper_6_io_in = swap;
  assign RetimeWrapper_6_clock = clock;
  assign RetimeWrapper_6_reset = reset;
  assign _T_61 = RetimeWrapper_6_io_out;
  assign RetimeWrapper_7_io_flow = 1'h1;
  assign RetimeWrapper_7_io_in = reset;
  assign RetimeWrapper_7_clock = clock;
  assign RetimeWrapper_7_reset = reset;
  assign _T_66 = RetimeWrapper_7_io_out;
  assign RetimeWrapper_8_io_flow = 1'h1;
  assign RetimeWrapper_8_io_in = swap;
  assign RetimeWrapper_8_clock = clock;
  assign RetimeWrapper_8_reset = reset;
  assign _T_70 = RetimeWrapper_8_io_out;
  assign RetimeWrapper_9_io_flow = 1'h1;
  assign RetimeWrapper_9_io_in = reset;
  assign RetimeWrapper_9_clock = clock;
  assign RetimeWrapper_9_reset = reset;
  assign _T_75 = RetimeWrapper_9_io_out;
  assign RetimeWrapper_10_io_flow = 1'h1;
  assign RetimeWrapper_10_io_in = _T_79;
  assign RetimeWrapper_10_clock = clock;
  assign RetimeWrapper_10_reset = reset;
  assign _T_83 = RetimeWrapper_10_io_out;
  assign RetimeWrapper_11_io_flow = 1'h1;
  assign RetimeWrapper_11_io_in = swap;
  assign RetimeWrapper_11_clock = clock;
  assign RetimeWrapper_11_reset = reset;
  assign _T_89 = RetimeWrapper_11_io_out;
  assign RetimeWrapper_12_io_flow = 1'h1;
  assign RetimeWrapper_12_io_in = reset;
  assign RetimeWrapper_12_clock = clock;
  assign RetimeWrapper_12_reset = reset;
  assign _T_94 = RetimeWrapper_12_io_out;
  assign RetimeWrapper_13_io_flow = 1'h1;
  assign RetimeWrapper_13_io_in = swap;
  assign RetimeWrapper_13_clock = clock;
  assign RetimeWrapper_13_reset = reset;
  assign _T_98 = RetimeWrapper_13_io_out;
  assign RetimeWrapper_14_io_flow = 1'h1;
  assign RetimeWrapper_14_io_in = reset;
  assign RetimeWrapper_14_clock = clock;
  assign RetimeWrapper_14_reset = reset;
  assign _T_103 = RetimeWrapper_14_io_out;
  assign RetimeWrapper_15_io_flow = 1'h1;
  assign RetimeWrapper_15_io_in = _T_107;
  assign RetimeWrapper_15_clock = clock;
  assign RetimeWrapper_15_reset = reset;
  assign _T_111 = RetimeWrapper_15_io_out;
  assign RetimeWrapper_16_io_flow = 1'h1;
  assign RetimeWrapper_16_io_in = swap;
  assign RetimeWrapper_16_clock = clock;
  assign RetimeWrapper_16_reset = reset;
  assign _T_117 = RetimeWrapper_16_io_out;
  assign RetimeWrapper_17_io_flow = 1'h1;
  assign RetimeWrapper_17_io_in = reset;
  assign RetimeWrapper_17_clock = clock;
  assign RetimeWrapper_17_reset = reset;
  assign _T_122 = RetimeWrapper_17_io_out;
  assign RetimeWrapper_18_io_flow = 1'h1;
  assign RetimeWrapper_18_io_in = swap;
  assign RetimeWrapper_18_clock = clock;
  assign RetimeWrapper_18_reset = reset;
  assign _T_126 = RetimeWrapper_18_io_out;
  assign RetimeWrapper_19_io_flow = 1'h1;
  assign RetimeWrapper_19_io_in = reset;
  assign RetimeWrapper_19_clock = clock;
  assign RetimeWrapper_19_reset = reset;
  assign _T_131 = RetimeWrapper_19_io_out;
  assign RetimeWrapper_20_io_flow = 1'h1;
  assign RetimeWrapper_20_io_in = _T_135;
  assign RetimeWrapper_20_clock = clock;
  assign RetimeWrapper_20_reset = reset;
  assign _T_139 = RetimeWrapper_20_io_out;
  assign RetimeWrapper_21_io_flow = 1'h1;
  assign RetimeWrapper_21_io_in = swap;
  assign RetimeWrapper_21_clock = clock;
  assign RetimeWrapper_21_reset = reset;
  assign _T_145 = RetimeWrapper_21_io_out;
  assign RetimeWrapper_22_io_flow = 1'h1;
  assign RetimeWrapper_22_io_in = reset;
  assign RetimeWrapper_22_clock = clock;
  assign RetimeWrapper_22_reset = reset;
  assign _T_150 = RetimeWrapper_22_io_out;
  assign RetimeWrapper_23_io_flow = 1'h1;
  assign RetimeWrapper_23_io_in = swap;
  assign RetimeWrapper_23_clock = clock;
  assign RetimeWrapper_23_reset = reset;
  assign _T_154 = RetimeWrapper_23_io_out;
  assign RetimeWrapper_24_io_flow = 1'h1;
  assign RetimeWrapper_24_io_in = reset;
  assign RetimeWrapper_24_clock = clock;
  assign RetimeWrapper_24_reset = reset;
  assign _T_159 = RetimeWrapper_24_io_out;
  assign statesIn_0_io_input_enable = swap;
  assign statesIn_0_clock = clock;
  assign statesIn_0_reset = reset;
  assign statesOut_0_io_input_enable = swap;
  assign statesOut_0_clock = clock;
  assign statesOut_0_reset = reset;
  assign statesOut_1_io_input_enable = swap;
  assign statesOut_1_clock = clock;
  assign statesOut_1_reset = reset;
  assign statesOut_2_io_input_enable = swap;
  assign statesOut_2_clock = clock;
  assign statesOut_2_reset = reset;
  assign statesOut_3_io_input_enable = swap;
  assign statesOut_3_clock = clock;
  assign statesOut_3_reset = reset;
  assign statesOut_4_io_input_enable = swap;
  assign statesOut_4_clock = clock;
  assign statesOut_4_reset = reset;
  assign _T_197_data = io_input_0_data;
  assign _T_197_enable = _T_198;
  assign _T_197_reset = io_input_0_reset;
  assign _T_203_data = io_input_0_data;
  assign _T_203_enable = _T_204;
  assign _T_203_reset = io_input_0_reset;
  assign _T_209_data = io_input_0_data;
  assign _T_209_enable = _T_210;
  assign _T_209_reset = io_input_0_reset;
  assign _T_215_data = io_input_0_data;
  assign _T_215_enable = _T_216;
  assign _T_215_reset = io_input_0_reset;
  assign _T_221_data = io_input_0_data;
  assign _T_221_enable = _T_222;
  assign _T_221_reset = io_input_0_reset;
  assign _T_273_0 = ff_0_io_output_data;
  assign _T_273_1 = ff_1_io_output_data;
  assign _T_273_2 = ff_2_io_output_data;
  assign _T_273_3 = ff_3_io_output_data;
  assign _T_273_4 = ff_4_io_output_data;
  assign _T_297 = _T_295;
  assign _T_310_0 = ff_0_io_output_data;
  assign _T_310_1 = ff_1_io_output_data;
  assign _T_310_2 = ff_2_io_output_data;
  assign _T_310_3 = ff_3_io_output_data;
  assign _T_310_4 = ff_4_io_output_data;
  assign _T_334 = _T_332;
  assign _T_384_0 = ff_0_io_output_data;
  assign _T_384_1 = ff_1_io_output_data;
  assign _T_384_2 = ff_2_io_output_data;
  assign _T_384_3 = ff_3_io_output_data;
  assign _T_384_4 = ff_4_io_output_data;
  assign _T_408 = _T_406;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_181 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_181 <= 1'h0;
    end else begin
      _T_181 <= _T_178;
    end
  end
endmodule
module RetimeWrapper_106(
  input        clock,
  input        reset,
  input  [2:0] io_in,
  output [2:0] io_out
);
  wire [2:0] sr_out;
  wire [2:0] sr_in;
  wire  sr_flow;
  wire  sr_reset;
  wire  sr_clock;
  RetimeShiftRegister #(.WIDTH(3), .STAGES(1)) sr (
    .out(sr_out),
    .in(sr_in),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out;
  assign sr_in = io_in;
  assign sr_flow = 1'h1;
  assign sr_reset = reset;
  assign sr_clock = clock;
endmodule
module NBufCtr_12(
  input        clock,
  input        reset,
  input        io_input_enable,
  output [2:0] io_output_count
);
  wire [2:0] _T_8;
  wire [3:0] _T_9;
  wire [2:0] _T_10;
  wire  _T_12;
  wire [3:0] _T_16;
  wire [3:0] _T_17;
  wire [2:0] _T_18;
  wire [2:0] _T_21;
  wire  _T_23;
  wire [3:0] _T_26;
  wire [3:0] _T_27;
  wire [2:0] _T_28;
  wire [2:0] _T_29;
  wire [2:0] _T_30;
  wire [2:0] _T_54;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire [2:0] RetimeWrapper_io_in;
  wire [2:0] RetimeWrapper_io_out;
  wire [2:0] _T_58;
  RetimeWrapper_106 RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_9 = _T_8 + 3'h0;
  assign _T_10 = _T_9[2:0];
  assign _T_12 = _T_10 >= 3'h4;
  assign _T_16 = _T_10 - 3'h4;
  assign _T_17 = $unsigned(_T_16);
  assign _T_18 = _T_17[2:0];
  assign _T_21 = _T_12 ? _T_18 : _T_10;
  assign _T_23 = _T_8 == 3'h0;
  assign _T_26 = _T_8 - 3'h1;
  assign _T_27 = $unsigned(_T_26);
  assign _T_28 = _T_27[2:0];
  assign _T_29 = _T_23 ? 3'h3 : _T_28;
  assign _T_30 = io_input_enable ? _T_29 : _T_8;
  assign _T_54 = reset ? 3'h0 : _T_30;
  assign io_output_count = _T_21;
  assign _T_8 = _T_58;
  assign RetimeWrapper_io_in = _T_54;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_58 = RetimeWrapper_io_out;
endmodule
module NBufCtr_13(
  input   clock,
  input   reset,
  input   io_input_enable
);
  wire [2:0] _T_8;
  wire  _T_25;
  wire [3:0] _T_28;
  wire [3:0] _T_29;
  wire [2:0] _T_30;
  wire [2:0] _T_31;
  wire [2:0] _T_32;
  wire [2:0] _T_55;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire [2:0] RetimeWrapper_io_in;
  wire [2:0] RetimeWrapper_io_out;
  wire [2:0] _T_59;
  RetimeWrapper_106 RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_25 = _T_8 == 3'h0;
  assign _T_28 = _T_8 - 3'h1;
  assign _T_29 = $unsigned(_T_28);
  assign _T_30 = _T_29[2:0];
  assign _T_31 = _T_25 ? 3'h3 : _T_30;
  assign _T_32 = io_input_enable ? _T_31 : _T_8;
  assign _T_55 = reset ? 3'h0 : _T_32;
  assign _T_8 = _T_59;
  assign RetimeWrapper_io_in = _T_55;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_59 = RetimeWrapper_io_out;
endmodule
module NBufCtr_14(
  input        clock,
  input        reset,
  input        io_input_enable,
  output [2:0] io_output_count
);
  wire [2:0] _T_8;
  wire [3:0] _T_10;
  wire [2:0] _T_11;
  wire  _T_13;
  wire [2:0] _T_14;
  wire [3:0] _T_16;
  wire [2:0] _T_17;
  wire [2:0] _T_18;
  wire [2:0] _T_19;
  wire [2:0] _T_23;
  wire  _T_25;
  wire [3:0] _T_28;
  wire [3:0] _T_29;
  wire [2:0] _T_30;
  wire [2:0] _T_31;
  wire [2:0] _T_32;
  wire [2:0] _T_55;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire [2:0] RetimeWrapper_io_in;
  wire [2:0] RetimeWrapper_io_out;
  wire [2:0] _T_59;
  RetimeWrapper_106 RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_10 = _T_8 + 3'h1;
  assign _T_11 = _T_10[2:0];
  assign _T_13 = _T_11 >= 3'h4;
  assign _T_14 = $signed(_T_8);
  assign _T_16 = $signed(_T_14) + $signed(-3'sh3);
  assign _T_17 = _T_16[2:0];
  assign _T_18 = $signed(_T_17);
  assign _T_19 = $unsigned(_T_18);
  assign _T_23 = _T_13 ? _T_19 : _T_11;
  assign _T_25 = _T_8 == 3'h0;
  assign _T_28 = _T_8 - 3'h1;
  assign _T_29 = $unsigned(_T_28);
  assign _T_30 = _T_29[2:0];
  assign _T_31 = _T_25 ? 3'h3 : _T_30;
  assign _T_32 = io_input_enable ? _T_31 : _T_8;
  assign _T_55 = reset ? 3'h0 : _T_32;
  assign io_output_count = _T_23;
  assign _T_8 = _T_59;
  assign RetimeWrapper_io_in = _T_55;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_59 = RetimeWrapper_io_out;
endmodule
module NBufCtr_15(
  input        clock,
  input        reset,
  input        io_input_enable,
  output [2:0] io_output_count
);
  wire [2:0] _T_8;
  wire [3:0] _T_10;
  wire [2:0] _T_11;
  wire  _T_13;
  wire [2:0] _T_14;
  wire [3:0] _T_16;
  wire [2:0] _T_17;
  wire [2:0] _T_18;
  wire [2:0] _T_19;
  wire [2:0] _T_23;
  wire  _T_25;
  wire [3:0] _T_28;
  wire [3:0] _T_29;
  wire [2:0] _T_30;
  wire [2:0] _T_31;
  wire [2:0] _T_32;
  wire [2:0] _T_55;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire [2:0] RetimeWrapper_io_in;
  wire [2:0] RetimeWrapper_io_out;
  wire [2:0] _T_59;
  RetimeWrapper_106 RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_10 = _T_8 + 3'h2;
  assign _T_11 = _T_10[2:0];
  assign _T_13 = _T_11 >= 3'h4;
  assign _T_14 = $signed(_T_8);
  assign _T_16 = $signed(_T_14) + $signed(-3'sh2);
  assign _T_17 = _T_16[2:0];
  assign _T_18 = $signed(_T_17);
  assign _T_19 = $unsigned(_T_18);
  assign _T_23 = _T_13 ? _T_19 : _T_11;
  assign _T_25 = _T_8 == 3'h0;
  assign _T_28 = _T_8 - 3'h1;
  assign _T_29 = $unsigned(_T_28);
  assign _T_30 = _T_29[2:0];
  assign _T_31 = _T_25 ? 3'h3 : _T_30;
  assign _T_32 = io_input_enable ? _T_31 : _T_8;
  assign _T_55 = reset ? 3'h0 : _T_32;
  assign io_output_count = _T_23;
  assign _T_8 = _T_59;
  assign RetimeWrapper_io_in = _T_55;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_59 = RetimeWrapper_io_out;
endmodule
module NBufCtr_16(
  input        clock,
  input        reset,
  input        io_input_enable,
  output [2:0] io_output_count
);
  wire [2:0] _T_8;
  wire [3:0] _T_10;
  wire [2:0] _T_11;
  wire  _T_13;
  wire [2:0] _T_14;
  wire [3:0] _T_16;
  wire [2:0] _T_17;
  wire [2:0] _T_18;
  wire [2:0] _T_19;
  wire [2:0] _T_23;
  wire  _T_25;
  wire [3:0] _T_28;
  wire [3:0] _T_29;
  wire [2:0] _T_30;
  wire [2:0] _T_31;
  wire [2:0] _T_32;
  wire [2:0] _T_55;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire [2:0] RetimeWrapper_io_in;
  wire [2:0] RetimeWrapper_io_out;
  wire [2:0] _T_59;
  RetimeWrapper_106 RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_10 = _T_8 + 3'h3;
  assign _T_11 = _T_10[2:0];
  assign _T_13 = _T_11 >= 3'h4;
  assign _T_14 = $signed(_T_8);
  assign _T_16 = $signed(_T_14) + $signed(-3'sh1);
  assign _T_17 = _T_16[2:0];
  assign _T_18 = $signed(_T_17);
  assign _T_19 = $unsigned(_T_18);
  assign _T_23 = _T_13 ? _T_19 : _T_11;
  assign _T_25 = _T_8 == 3'h0;
  assign _T_28 = _T_8 - 3'h1;
  assign _T_29 = $unsigned(_T_28);
  assign _T_30 = _T_29[2:0];
  assign _T_31 = _T_25 ? 3'h3 : _T_30;
  assign _T_32 = io_input_enable ? _T_31 : _T_8;
  assign _T_55 = reset ? 3'h0 : _T_32;
  assign io_output_count = _T_23;
  assign _T_8 = _T_59;
  assign RetimeWrapper_io_in = _T_55;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_59 = RetimeWrapper_io_out;
endmodule
module NBufFF_2(
  input         clock,
  input         reset,
  input         io_sEn_0,
  input         io_sEn_1,
  input         io_sEn_2,
  input         io_sEn_3,
  input         io_sDone_0,
  input         io_sDone_1,
  input         io_sDone_2,
  input         io_sDone_3,
  input  [31:0] io_input_0_data,
  input         io_input_0_enable,
  input         io_input_0_reset,
  output [31:0] io_output_1_data,
  output [31:0] io_output_2_data,
  output [31:0] io_output_3_data
);
  wire  ff_0_clock;
  wire  ff_0_reset;
  wire [31:0] ff_0_io_input_0_data;
  wire [31:0] ff_0_io_input_0_init;
  wire  ff_0_io_input_0_enable;
  wire  ff_0_io_input_0_reset;
  wire [31:0] ff_0_io_output_data;
  wire  ff_1_clock;
  wire  ff_1_reset;
  wire [31:0] ff_1_io_input_0_data;
  wire [31:0] ff_1_io_input_0_init;
  wire  ff_1_io_input_0_enable;
  wire  ff_1_io_input_0_reset;
  wire [31:0] ff_1_io_output_data;
  wire  ff_2_clock;
  wire  ff_2_reset;
  wire [31:0] ff_2_io_input_0_data;
  wire [31:0] ff_2_io_input_0_init;
  wire  ff_2_io_input_0_enable;
  wire  ff_2_io_input_0_reset;
  wire [31:0] ff_2_io_output_data;
  wire  ff_3_clock;
  wire  ff_3_reset;
  wire [31:0] ff_3_io_input_0_data;
  wire [31:0] ff_3_io_input_0_init;
  wire  ff_3_io_input_0_enable;
  wire  ff_3_io_input_0_reset;
  wire [31:0] ff_3_io_output_data;
  wire  sEn_latch_0_clock;
  wire  sEn_latch_0_reset;
  wire  sEn_latch_0_io_input_set;
  wire  sEn_latch_0_io_input_reset;
  wire  sEn_latch_0_io_input_asyn_reset;
  wire  sEn_latch_0_io_output_data;
  wire  sEn_latch_1_clock;
  wire  sEn_latch_1_reset;
  wire  sEn_latch_1_io_input_set;
  wire  sEn_latch_1_io_input_reset;
  wire  sEn_latch_1_io_input_asyn_reset;
  wire  sEn_latch_1_io_output_data;
  wire  sEn_latch_2_clock;
  wire  sEn_latch_2_reset;
  wire  sEn_latch_2_io_input_set;
  wire  sEn_latch_2_io_input_reset;
  wire  sEn_latch_2_io_input_asyn_reset;
  wire  sEn_latch_2_io_output_data;
  wire  sEn_latch_3_clock;
  wire  sEn_latch_3_reset;
  wire  sEn_latch_3_io_input_set;
  wire  sEn_latch_3_io_input_reset;
  wire  sEn_latch_3_io_input_asyn_reset;
  wire  sEn_latch_3_io_output_data;
  wire  sDone_latch_0_clock;
  wire  sDone_latch_0_reset;
  wire  sDone_latch_0_io_input_set;
  wire  sDone_latch_0_io_input_reset;
  wire  sDone_latch_0_io_input_asyn_reset;
  wire  sDone_latch_0_io_output_data;
  wire  sDone_latch_1_clock;
  wire  sDone_latch_1_reset;
  wire  sDone_latch_1_io_input_set;
  wire  sDone_latch_1_io_input_reset;
  wire  sDone_latch_1_io_input_asyn_reset;
  wire  sDone_latch_1_io_output_data;
  wire  sDone_latch_2_clock;
  wire  sDone_latch_2_reset;
  wire  sDone_latch_2_io_input_set;
  wire  sDone_latch_2_io_input_reset;
  wire  sDone_latch_2_io_input_asyn_reset;
  wire  sDone_latch_2_io_output_data;
  wire  sDone_latch_3_clock;
  wire  sDone_latch_3_reset;
  wire  sDone_latch_3_io_input_set;
  wire  sDone_latch_3_io_input_reset;
  wire  sDone_latch_3_io_input_asyn_reset;
  wire  sDone_latch_3_io_output_data;
  wire  swap;
  wire  _T_20;
  wire  _T_21;
  wire  _T_22;
  wire  _T_23;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire  RetimeWrapper_io_flow;
  wire  RetimeWrapper_io_in;
  wire  RetimeWrapper_io_out;
  wire  _T_27;
  wire  _T_28;
  wire  _T_29;
  wire  RetimeWrapper_1_clock;
  wire  RetimeWrapper_1_reset;
  wire  RetimeWrapper_1_io_flow;
  wire  RetimeWrapper_1_io_in;
  wire  RetimeWrapper_1_io_out;
  wire  _T_33;
  wire  _T_34;
  wire  RetimeWrapper_2_clock;
  wire  RetimeWrapper_2_reset;
  wire  RetimeWrapper_2_io_flow;
  wire  RetimeWrapper_2_io_in;
  wire  RetimeWrapper_2_io_out;
  wire  _T_38;
  wire  RetimeWrapper_3_clock;
  wire  RetimeWrapper_3_reset;
  wire  RetimeWrapper_3_io_flow;
  wire  RetimeWrapper_3_io_in;
  wire  RetimeWrapper_3_io_out;
  wire  _T_42;
  wire  _T_43;
  wire  RetimeWrapper_4_clock;
  wire  RetimeWrapper_4_reset;
  wire  RetimeWrapper_4_io_flow;
  wire  RetimeWrapper_4_io_in;
  wire  RetimeWrapper_4_io_out;
  wire  _T_47;
  wire  _T_48;
  wire  _T_49;
  wire  _T_50;
  wire  _T_51;
  wire  RetimeWrapper_5_clock;
  wire  RetimeWrapper_5_reset;
  wire  RetimeWrapper_5_io_flow;
  wire  RetimeWrapper_5_io_in;
  wire  RetimeWrapper_5_io_out;
  wire  _T_55;
  wire  _T_56;
  wire  _T_57;
  wire  RetimeWrapper_6_clock;
  wire  RetimeWrapper_6_reset;
  wire  RetimeWrapper_6_io_flow;
  wire  RetimeWrapper_6_io_in;
  wire  RetimeWrapper_6_io_out;
  wire  _T_61;
  wire  _T_62;
  wire  RetimeWrapper_7_clock;
  wire  RetimeWrapper_7_reset;
  wire  RetimeWrapper_7_io_flow;
  wire  RetimeWrapper_7_io_in;
  wire  RetimeWrapper_7_io_out;
  wire  _T_66;
  wire  RetimeWrapper_8_clock;
  wire  RetimeWrapper_8_reset;
  wire  RetimeWrapper_8_io_flow;
  wire  RetimeWrapper_8_io_in;
  wire  RetimeWrapper_8_io_out;
  wire  _T_70;
  wire  _T_71;
  wire  RetimeWrapper_9_clock;
  wire  RetimeWrapper_9_reset;
  wire  RetimeWrapper_9_io_flow;
  wire  RetimeWrapper_9_io_in;
  wire  RetimeWrapper_9_io_out;
  wire  _T_75;
  wire  _T_76;
  wire  _T_77;
  wire  _T_78;
  wire  _T_79;
  wire  RetimeWrapper_10_clock;
  wire  RetimeWrapper_10_reset;
  wire  RetimeWrapper_10_io_flow;
  wire  RetimeWrapper_10_io_in;
  wire  RetimeWrapper_10_io_out;
  wire  _T_83;
  wire  _T_84;
  wire  _T_85;
  wire  RetimeWrapper_11_clock;
  wire  RetimeWrapper_11_reset;
  wire  RetimeWrapper_11_io_flow;
  wire  RetimeWrapper_11_io_in;
  wire  RetimeWrapper_11_io_out;
  wire  _T_89;
  wire  _T_90;
  wire  RetimeWrapper_12_clock;
  wire  RetimeWrapper_12_reset;
  wire  RetimeWrapper_12_io_flow;
  wire  RetimeWrapper_12_io_in;
  wire  RetimeWrapper_12_io_out;
  wire  _T_94;
  wire  RetimeWrapper_13_clock;
  wire  RetimeWrapper_13_reset;
  wire  RetimeWrapper_13_io_flow;
  wire  RetimeWrapper_13_io_in;
  wire  RetimeWrapper_13_io_out;
  wire  _T_98;
  wire  _T_99;
  wire  RetimeWrapper_14_clock;
  wire  RetimeWrapper_14_reset;
  wire  RetimeWrapper_14_io_flow;
  wire  RetimeWrapper_14_io_in;
  wire  RetimeWrapper_14_io_out;
  wire  _T_103;
  wire  _T_104;
  wire  _T_105;
  wire  _T_106;
  wire  _T_107;
  wire  RetimeWrapper_15_clock;
  wire  RetimeWrapper_15_reset;
  wire  RetimeWrapper_15_io_flow;
  wire  RetimeWrapper_15_io_in;
  wire  RetimeWrapper_15_io_out;
  wire  _T_111;
  wire  _T_112;
  wire  _T_113;
  wire  RetimeWrapper_16_clock;
  wire  RetimeWrapper_16_reset;
  wire  RetimeWrapper_16_io_flow;
  wire  RetimeWrapper_16_io_in;
  wire  RetimeWrapper_16_io_out;
  wire  _T_117;
  wire  _T_118;
  wire  RetimeWrapper_17_clock;
  wire  RetimeWrapper_17_reset;
  wire  RetimeWrapper_17_io_flow;
  wire  RetimeWrapper_17_io_in;
  wire  RetimeWrapper_17_io_out;
  wire  _T_122;
  wire  RetimeWrapper_18_clock;
  wire  RetimeWrapper_18_reset;
  wire  RetimeWrapper_18_io_flow;
  wire  RetimeWrapper_18_io_in;
  wire  RetimeWrapper_18_io_out;
  wire  _T_126;
  wire  _T_127;
  wire  RetimeWrapper_19_clock;
  wire  RetimeWrapper_19_reset;
  wire  RetimeWrapper_19_io_flow;
  wire  RetimeWrapper_19_io_in;
  wire  RetimeWrapper_19_io_out;
  wire  _T_131;
  wire  _T_132;
  wire  _T_133;
  wire  anyEnabled;
  wire  _T_134;
  wire  _T_135;
  wire  _T_136;
  wire  _T_137;
  wire  _T_138;
  wire  _T_139;
  wire  _T_140;
  wire  _T_141;
  wire  _T_142;
  wire  _T_143;
  wire  _T_144;
  wire  _T_145;
  wire  _T_146;
  reg  _T_149;
  reg [31:0] _RAND_0;
  wire  _T_155;
  wire  statesIn_0_clock;
  wire  statesIn_0_reset;
  wire  statesIn_0_io_input_enable;
  wire [2:0] statesIn_0_io_output_count;
  wire  statesOut_0_clock;
  wire  statesOut_0_reset;
  wire  statesOut_0_io_input_enable;
  wire  statesOut_1_clock;
  wire  statesOut_1_reset;
  wire  statesOut_1_io_input_enable;
  wire [2:0] statesOut_1_io_output_count;
  wire  statesOut_2_clock;
  wire  statesOut_2_reset;
  wire  statesOut_2_io_input_enable;
  wire [2:0] statesOut_2_io_output_count;
  wire  statesOut_3_clock;
  wire  statesOut_3_reset;
  wire  statesOut_3_io_input_enable;
  wire [2:0] statesOut_3_io_output_count;
  wire  _T_162;
  wire [31:0] _T_164_data;
  wire  _T_164_enable;
  wire  _T_164_reset;
  wire  _T_165;
  wire  _T_168;
  wire [31:0] _T_170_data;
  wire  _T_170_enable;
  wire  _T_170_reset;
  wire  _T_171;
  wire  _T_174;
  wire [31:0] _T_176_data;
  wire  _T_176_enable;
  wire  _T_176_reset;
  wire  _T_177;
  wire  _T_180;
  wire [31:0] _T_182_data;
  wire  _T_182_enable;
  wire  _T_182_reset;
  wire  _T_183;
  wire  _T_217;
  wire  _T_219;
  wire  _T_221;
  wire  _T_223;
  wire [31:0] _T_226_0;
  wire [31:0] _T_226_1;
  wire [31:0] _T_226_2;
  wire [31:0] _T_226_3;
  wire [31:0] _T_235;
  wire [31:0] _T_237;
  wire [31:0] _T_239;
  wire [31:0] _T_241;
  wire [31:0] _T_242;
  wire [31:0] _T_243;
  wire [31:0] _T_244;
  wire [31:0] _T_246;
  wire  _T_248;
  wire  _T_250;
  wire  _T_252;
  wire  _T_254;
  wire [31:0] _T_257_0;
  wire [31:0] _T_257_1;
  wire [31:0] _T_257_2;
  wire [31:0] _T_257_3;
  wire [31:0] _T_266;
  wire [31:0] _T_268;
  wire [31:0] _T_270;
  wire [31:0] _T_272;
  wire [31:0] _T_273;
  wire [31:0] _T_274;
  wire [31:0] _T_275;
  wire [31:0] _T_277;
  wire  _T_279;
  wire  _T_281;
  wire  _T_283;
  wire  _T_285;
  wire [31:0] _T_288_0;
  wire [31:0] _T_288_1;
  wire [31:0] _T_288_2;
  wire [31:0] _T_288_3;
  wire [31:0] _T_297;
  wire [31:0] _T_299;
  wire [31:0] _T_301;
  wire [31:0] _T_303;
  wire [31:0] _T_304;
  wire [31:0] _T_305;
  wire [31:0] _T_306;
  wire [31:0] _T_308;
  FF_1 ff_0 (
    .clock(ff_0_clock),
    .reset(ff_0_reset),
    .io_input_0_data(ff_0_io_input_0_data),
    .io_input_0_init(ff_0_io_input_0_init),
    .io_input_0_enable(ff_0_io_input_0_enable),
    .io_input_0_reset(ff_0_io_input_0_reset),
    .io_output_data(ff_0_io_output_data)
  );
  FF_1 ff_1 (
    .clock(ff_1_clock),
    .reset(ff_1_reset),
    .io_input_0_data(ff_1_io_input_0_data),
    .io_input_0_init(ff_1_io_input_0_init),
    .io_input_0_enable(ff_1_io_input_0_enable),
    .io_input_0_reset(ff_1_io_input_0_reset),
    .io_output_data(ff_1_io_output_data)
  );
  FF_1 ff_2 (
    .clock(ff_2_clock),
    .reset(ff_2_reset),
    .io_input_0_data(ff_2_io_input_0_data),
    .io_input_0_init(ff_2_io_input_0_init),
    .io_input_0_enable(ff_2_io_input_0_enable),
    .io_input_0_reset(ff_2_io_input_0_reset),
    .io_output_data(ff_2_io_output_data)
  );
  FF_1 ff_3 (
    .clock(ff_3_clock),
    .reset(ff_3_reset),
    .io_input_0_data(ff_3_io_input_0_data),
    .io_input_0_init(ff_3_io_input_0_init),
    .io_input_0_enable(ff_3_io_input_0_enable),
    .io_input_0_reset(ff_3_io_input_0_reset),
    .io_output_data(ff_3_io_output_data)
  );
  SRFF sEn_latch_0 (
    .clock(sEn_latch_0_clock),
    .reset(sEn_latch_0_reset),
    .io_input_set(sEn_latch_0_io_input_set),
    .io_input_reset(sEn_latch_0_io_input_reset),
    .io_input_asyn_reset(sEn_latch_0_io_input_asyn_reset),
    .io_output_data(sEn_latch_0_io_output_data)
  );
  SRFF sEn_latch_1 (
    .clock(sEn_latch_1_clock),
    .reset(sEn_latch_1_reset),
    .io_input_set(sEn_latch_1_io_input_set),
    .io_input_reset(sEn_latch_1_io_input_reset),
    .io_input_asyn_reset(sEn_latch_1_io_input_asyn_reset),
    .io_output_data(sEn_latch_1_io_output_data)
  );
  SRFF sEn_latch_2 (
    .clock(sEn_latch_2_clock),
    .reset(sEn_latch_2_reset),
    .io_input_set(sEn_latch_2_io_input_set),
    .io_input_reset(sEn_latch_2_io_input_reset),
    .io_input_asyn_reset(sEn_latch_2_io_input_asyn_reset),
    .io_output_data(sEn_latch_2_io_output_data)
  );
  SRFF sEn_latch_3 (
    .clock(sEn_latch_3_clock),
    .reset(sEn_latch_3_reset),
    .io_input_set(sEn_latch_3_io_input_set),
    .io_input_reset(sEn_latch_3_io_input_reset),
    .io_input_asyn_reset(sEn_latch_3_io_input_asyn_reset),
    .io_output_data(sEn_latch_3_io_output_data)
  );
  SRFF sDone_latch_0 (
    .clock(sDone_latch_0_clock),
    .reset(sDone_latch_0_reset),
    .io_input_set(sDone_latch_0_io_input_set),
    .io_input_reset(sDone_latch_0_io_input_reset),
    .io_input_asyn_reset(sDone_latch_0_io_input_asyn_reset),
    .io_output_data(sDone_latch_0_io_output_data)
  );
  SRFF sDone_latch_1 (
    .clock(sDone_latch_1_clock),
    .reset(sDone_latch_1_reset),
    .io_input_set(sDone_latch_1_io_input_set),
    .io_input_reset(sDone_latch_1_io_input_reset),
    .io_input_asyn_reset(sDone_latch_1_io_input_asyn_reset),
    .io_output_data(sDone_latch_1_io_output_data)
  );
  SRFF sDone_latch_2 (
    .clock(sDone_latch_2_clock),
    .reset(sDone_latch_2_reset),
    .io_input_set(sDone_latch_2_io_input_set),
    .io_input_reset(sDone_latch_2_io_input_reset),
    .io_input_asyn_reset(sDone_latch_2_io_input_asyn_reset),
    .io_output_data(sDone_latch_2_io_output_data)
  );
  SRFF sDone_latch_3 (
    .clock(sDone_latch_3_clock),
    .reset(sDone_latch_3_reset),
    .io_input_set(sDone_latch_3_io_input_set),
    .io_input_reset(sDone_latch_3_io_input_reset),
    .io_input_asyn_reset(sDone_latch_3_io_input_asyn_reset),
    .io_output_data(sDone_latch_3_io_output_data)
  );
  RetimeWrapper RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 (
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 (
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 (
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 (
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 (
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 (
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 (
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper RetimeWrapper_8 (
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper RetimeWrapper_9 (
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper RetimeWrapper_10 (
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper RetimeWrapper_11 (
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper RetimeWrapper_12 (
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper RetimeWrapper_13 (
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper RetimeWrapper_14 (
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper RetimeWrapper_15 (
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper RetimeWrapper_16 (
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper RetimeWrapper_17 (
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper RetimeWrapper_18 (
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper RetimeWrapper_19 (
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  NBufCtr_12 statesIn_0 (
    .clock(statesIn_0_clock),
    .reset(statesIn_0_reset),
    .io_input_enable(statesIn_0_io_input_enable),
    .io_output_count(statesIn_0_io_output_count)
  );
  NBufCtr_13 statesOut_0 (
    .clock(statesOut_0_clock),
    .reset(statesOut_0_reset),
    .io_input_enable(statesOut_0_io_input_enable)
  );
  NBufCtr_14 statesOut_1 (
    .clock(statesOut_1_clock),
    .reset(statesOut_1_reset),
    .io_input_enable(statesOut_1_io_input_enable),
    .io_output_count(statesOut_1_io_output_count)
  );
  NBufCtr_15 statesOut_2 (
    .clock(statesOut_2_clock),
    .reset(statesOut_2_reset),
    .io_input_enable(statesOut_2_io_input_enable),
    .io_output_count(statesOut_2_io_output_count)
  );
  NBufCtr_16 statesOut_3 (
    .clock(statesOut_3_clock),
    .reset(statesOut_3_reset),
    .io_input_enable(statesOut_3_io_input_enable),
    .io_output_count(statesOut_3_io_output_count)
  );
  assign _T_20 = ~ io_sDone_0;
  assign _T_21 = io_sEn_0 & _T_20;
  assign _T_22 = io_sEn_0 & io_sDone_0;
  assign _T_23 = ~ io_sEn_0;
  assign _T_28 = _T_22 & _T_27;
  assign _T_29 = _T_21 | _T_28;
  assign _T_34 = swap | _T_33;
  assign _T_43 = swap | _T_42;
  assign _T_48 = ~ io_sDone_1;
  assign _T_49 = io_sEn_1 & _T_48;
  assign _T_50 = io_sEn_1 & io_sDone_1;
  assign _T_51 = ~ io_sEn_1;
  assign _T_56 = _T_50 & _T_55;
  assign _T_57 = _T_49 | _T_56;
  assign _T_62 = swap | _T_61;
  assign _T_71 = swap | _T_70;
  assign _T_76 = ~ io_sDone_2;
  assign _T_77 = io_sEn_2 & _T_76;
  assign _T_78 = io_sEn_2 & io_sDone_2;
  assign _T_79 = ~ io_sEn_2;
  assign _T_84 = _T_78 & _T_83;
  assign _T_85 = _T_77 | _T_84;
  assign _T_90 = swap | _T_89;
  assign _T_99 = swap | _T_98;
  assign _T_104 = ~ io_sDone_3;
  assign _T_105 = io_sEn_3 & _T_104;
  assign _T_106 = io_sEn_3 & io_sDone_3;
  assign _T_107 = ~ io_sEn_3;
  assign _T_112 = _T_106 & _T_111;
  assign _T_113 = _T_105 | _T_112;
  assign _T_118 = swap | _T_117;
  assign _T_127 = swap | _T_126;
  assign _T_132 = sEn_latch_0_io_output_data | sEn_latch_1_io_output_data;
  assign _T_133 = _T_132 | sEn_latch_2_io_output_data;
  assign anyEnabled = _T_133 | sEn_latch_3_io_output_data;
  assign _T_134 = sDone_latch_0_io_output_data | io_sDone_0;
  assign _T_135 = sEn_latch_0_io_output_data == _T_134;
  assign _T_136 = sDone_latch_1_io_output_data | io_sDone_1;
  assign _T_137 = sEn_latch_1_io_output_data == _T_136;
  assign _T_138 = sDone_latch_2_io_output_data | io_sDone_2;
  assign _T_139 = sEn_latch_2_io_output_data == _T_138;
  assign _T_140 = sDone_latch_3_io_output_data | io_sDone_3;
  assign _T_141 = sEn_latch_3_io_output_data == _T_140;
  assign _T_142 = _T_135 & _T_137;
  assign _T_143 = _T_142 & _T_139;
  assign _T_144 = _T_143 & _T_141;
  assign _T_145 = _T_144 & anyEnabled;
  assign _T_146 = ~ _T_145;
  assign _T_155 = _T_145 & _T_149;
  assign _T_162 = statesIn_0_io_output_count == 3'h0;
  assign _T_165 = io_input_0_enable & _T_162;
  assign _T_168 = statesIn_0_io_output_count == 3'h1;
  assign _T_171 = io_input_0_enable & _T_168;
  assign _T_174 = statesIn_0_io_output_count == 3'h2;
  assign _T_177 = io_input_0_enable & _T_174;
  assign _T_180 = statesIn_0_io_output_count == 3'h3;
  assign _T_183 = io_input_0_enable & _T_180;
  assign _T_217 = statesOut_1_io_output_count == 3'h0;
  assign _T_219 = statesOut_1_io_output_count == 3'h1;
  assign _T_221 = statesOut_1_io_output_count == 3'h2;
  assign _T_223 = statesOut_1_io_output_count == 3'h3;
  assign _T_235 = _T_217 ? _T_226_0 : 32'h0;
  assign _T_237 = _T_219 ? _T_226_1 : 32'h0;
  assign _T_239 = _T_221 ? _T_226_2 : 32'h0;
  assign _T_241 = _T_223 ? _T_226_3 : 32'h0;
  assign _T_242 = _T_235 | _T_237;
  assign _T_243 = _T_242 | _T_239;
  assign _T_244 = _T_243 | _T_241;
  assign _T_248 = statesOut_2_io_output_count == 3'h0;
  assign _T_250 = statesOut_2_io_output_count == 3'h1;
  assign _T_252 = statesOut_2_io_output_count == 3'h2;
  assign _T_254 = statesOut_2_io_output_count == 3'h3;
  assign _T_266 = _T_248 ? _T_257_0 : 32'h0;
  assign _T_268 = _T_250 ? _T_257_1 : 32'h0;
  assign _T_270 = _T_252 ? _T_257_2 : 32'h0;
  assign _T_272 = _T_254 ? _T_257_3 : 32'h0;
  assign _T_273 = _T_266 | _T_268;
  assign _T_274 = _T_273 | _T_270;
  assign _T_275 = _T_274 | _T_272;
  assign _T_279 = statesOut_3_io_output_count == 3'h0;
  assign _T_281 = statesOut_3_io_output_count == 3'h1;
  assign _T_283 = statesOut_3_io_output_count == 3'h2;
  assign _T_285 = statesOut_3_io_output_count == 3'h3;
  assign _T_297 = _T_279 ? _T_288_0 : 32'h0;
  assign _T_299 = _T_281 ? _T_288_1 : 32'h0;
  assign _T_301 = _T_283 ? _T_288_2 : 32'h0;
  assign _T_303 = _T_285 ? _T_288_3 : 32'h0;
  assign _T_304 = _T_297 | _T_299;
  assign _T_305 = _T_304 | _T_301;
  assign _T_306 = _T_305 | _T_303;
  assign io_output_1_data = _T_246;
  assign io_output_2_data = _T_277;
  assign io_output_3_data = _T_308;
  assign ff_0_io_input_0_data = _T_164_data;
  assign ff_0_io_input_0_init = 32'h0;
  assign ff_0_io_input_0_enable = _T_164_enable;
  assign ff_0_io_input_0_reset = _T_164_reset;
  assign ff_0_clock = clock;
  assign ff_0_reset = reset;
  assign ff_1_io_input_0_data = _T_170_data;
  assign ff_1_io_input_0_init = 32'h0;
  assign ff_1_io_input_0_enable = _T_170_enable;
  assign ff_1_io_input_0_reset = _T_170_reset;
  assign ff_1_clock = clock;
  assign ff_1_reset = reset;
  assign ff_2_io_input_0_data = _T_176_data;
  assign ff_2_io_input_0_init = 32'h0;
  assign ff_2_io_input_0_enable = _T_176_enable;
  assign ff_2_io_input_0_reset = _T_176_reset;
  assign ff_2_clock = clock;
  assign ff_2_reset = reset;
  assign ff_3_io_input_0_data = _T_182_data;
  assign ff_3_io_input_0_init = 32'h0;
  assign ff_3_io_input_0_enable = _T_182_enable;
  assign ff_3_io_input_0_reset = _T_182_reset;
  assign ff_3_clock = clock;
  assign ff_3_reset = reset;
  assign sEn_latch_0_io_input_set = _T_29;
  assign sEn_latch_0_io_input_reset = _T_34;
  assign sEn_latch_0_io_input_asyn_reset = _T_38;
  assign sEn_latch_0_clock = clock;
  assign sEn_latch_0_reset = reset;
  assign sEn_latch_1_io_input_set = _T_57;
  assign sEn_latch_1_io_input_reset = _T_62;
  assign sEn_latch_1_io_input_asyn_reset = _T_66;
  assign sEn_latch_1_clock = clock;
  assign sEn_latch_1_reset = reset;
  assign sEn_latch_2_io_input_set = _T_85;
  assign sEn_latch_2_io_input_reset = _T_90;
  assign sEn_latch_2_io_input_asyn_reset = _T_94;
  assign sEn_latch_2_clock = clock;
  assign sEn_latch_2_reset = reset;
  assign sEn_latch_3_io_input_set = _T_113;
  assign sEn_latch_3_io_input_reset = _T_118;
  assign sEn_latch_3_io_input_asyn_reset = _T_122;
  assign sEn_latch_3_clock = clock;
  assign sEn_latch_3_reset = reset;
  assign sDone_latch_0_io_input_set = io_sDone_0;
  assign sDone_latch_0_io_input_reset = _T_43;
  assign sDone_latch_0_io_input_asyn_reset = _T_47;
  assign sDone_latch_0_clock = clock;
  assign sDone_latch_0_reset = reset;
  assign sDone_latch_1_io_input_set = io_sDone_1;
  assign sDone_latch_1_io_input_reset = _T_71;
  assign sDone_latch_1_io_input_asyn_reset = _T_75;
  assign sDone_latch_1_clock = clock;
  assign sDone_latch_1_reset = reset;
  assign sDone_latch_2_io_input_set = io_sDone_2;
  assign sDone_latch_2_io_input_reset = _T_99;
  assign sDone_latch_2_io_input_asyn_reset = _T_103;
  assign sDone_latch_2_clock = clock;
  assign sDone_latch_2_reset = reset;
  assign sDone_latch_3_io_input_set = io_sDone_3;
  assign sDone_latch_3_io_input_reset = _T_127;
  assign sDone_latch_3_io_input_asyn_reset = _T_131;
  assign sDone_latch_3_clock = clock;
  assign sDone_latch_3_reset = reset;
  assign swap = _T_155;
  assign RetimeWrapper_io_flow = 1'h1;
  assign RetimeWrapper_io_in = _T_23;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_27 = RetimeWrapper_io_out;
  assign RetimeWrapper_1_io_flow = 1'h1;
  assign RetimeWrapper_1_io_in = swap;
  assign RetimeWrapper_1_clock = clock;
  assign RetimeWrapper_1_reset = reset;
  assign _T_33 = RetimeWrapper_1_io_out;
  assign RetimeWrapper_2_io_flow = 1'h1;
  assign RetimeWrapper_2_io_in = reset;
  assign RetimeWrapper_2_clock = clock;
  assign RetimeWrapper_2_reset = reset;
  assign _T_38 = RetimeWrapper_2_io_out;
  assign RetimeWrapper_3_io_flow = 1'h1;
  assign RetimeWrapper_3_io_in = swap;
  assign RetimeWrapper_3_clock = clock;
  assign RetimeWrapper_3_reset = reset;
  assign _T_42 = RetimeWrapper_3_io_out;
  assign RetimeWrapper_4_io_flow = 1'h1;
  assign RetimeWrapper_4_io_in = reset;
  assign RetimeWrapper_4_clock = clock;
  assign RetimeWrapper_4_reset = reset;
  assign _T_47 = RetimeWrapper_4_io_out;
  assign RetimeWrapper_5_io_flow = 1'h1;
  assign RetimeWrapper_5_io_in = _T_51;
  assign RetimeWrapper_5_clock = clock;
  assign RetimeWrapper_5_reset = reset;
  assign _T_55 = RetimeWrapper_5_io_out;
  assign RetimeWrapper_6_io_flow = 1'h1;
  assign RetimeWrapper_6_io_in = swap;
  assign RetimeWrapper_6_clock = clock;
  assign RetimeWrapper_6_reset = reset;
  assign _T_61 = RetimeWrapper_6_io_out;
  assign RetimeWrapper_7_io_flow = 1'h1;
  assign RetimeWrapper_7_io_in = reset;
  assign RetimeWrapper_7_clock = clock;
  assign RetimeWrapper_7_reset = reset;
  assign _T_66 = RetimeWrapper_7_io_out;
  assign RetimeWrapper_8_io_flow = 1'h1;
  assign RetimeWrapper_8_io_in = swap;
  assign RetimeWrapper_8_clock = clock;
  assign RetimeWrapper_8_reset = reset;
  assign _T_70 = RetimeWrapper_8_io_out;
  assign RetimeWrapper_9_io_flow = 1'h1;
  assign RetimeWrapper_9_io_in = reset;
  assign RetimeWrapper_9_clock = clock;
  assign RetimeWrapper_9_reset = reset;
  assign _T_75 = RetimeWrapper_9_io_out;
  assign RetimeWrapper_10_io_flow = 1'h1;
  assign RetimeWrapper_10_io_in = _T_79;
  assign RetimeWrapper_10_clock = clock;
  assign RetimeWrapper_10_reset = reset;
  assign _T_83 = RetimeWrapper_10_io_out;
  assign RetimeWrapper_11_io_flow = 1'h1;
  assign RetimeWrapper_11_io_in = swap;
  assign RetimeWrapper_11_clock = clock;
  assign RetimeWrapper_11_reset = reset;
  assign _T_89 = RetimeWrapper_11_io_out;
  assign RetimeWrapper_12_io_flow = 1'h1;
  assign RetimeWrapper_12_io_in = reset;
  assign RetimeWrapper_12_clock = clock;
  assign RetimeWrapper_12_reset = reset;
  assign _T_94 = RetimeWrapper_12_io_out;
  assign RetimeWrapper_13_io_flow = 1'h1;
  assign RetimeWrapper_13_io_in = swap;
  assign RetimeWrapper_13_clock = clock;
  assign RetimeWrapper_13_reset = reset;
  assign _T_98 = RetimeWrapper_13_io_out;
  assign RetimeWrapper_14_io_flow = 1'h1;
  assign RetimeWrapper_14_io_in = reset;
  assign RetimeWrapper_14_clock = clock;
  assign RetimeWrapper_14_reset = reset;
  assign _T_103 = RetimeWrapper_14_io_out;
  assign RetimeWrapper_15_io_flow = 1'h1;
  assign RetimeWrapper_15_io_in = _T_107;
  assign RetimeWrapper_15_clock = clock;
  assign RetimeWrapper_15_reset = reset;
  assign _T_111 = RetimeWrapper_15_io_out;
  assign RetimeWrapper_16_io_flow = 1'h1;
  assign RetimeWrapper_16_io_in = swap;
  assign RetimeWrapper_16_clock = clock;
  assign RetimeWrapper_16_reset = reset;
  assign _T_117 = RetimeWrapper_16_io_out;
  assign RetimeWrapper_17_io_flow = 1'h1;
  assign RetimeWrapper_17_io_in = reset;
  assign RetimeWrapper_17_clock = clock;
  assign RetimeWrapper_17_reset = reset;
  assign _T_122 = RetimeWrapper_17_io_out;
  assign RetimeWrapper_18_io_flow = 1'h1;
  assign RetimeWrapper_18_io_in = swap;
  assign RetimeWrapper_18_clock = clock;
  assign RetimeWrapper_18_reset = reset;
  assign _T_126 = RetimeWrapper_18_io_out;
  assign RetimeWrapper_19_io_flow = 1'h1;
  assign RetimeWrapper_19_io_in = reset;
  assign RetimeWrapper_19_clock = clock;
  assign RetimeWrapper_19_reset = reset;
  assign _T_131 = RetimeWrapper_19_io_out;
  assign statesIn_0_io_input_enable = swap;
  assign statesIn_0_clock = clock;
  assign statesIn_0_reset = reset;
  assign statesOut_0_io_input_enable = swap;
  assign statesOut_0_clock = clock;
  assign statesOut_0_reset = reset;
  assign statesOut_1_io_input_enable = swap;
  assign statesOut_1_clock = clock;
  assign statesOut_1_reset = reset;
  assign statesOut_2_io_input_enable = swap;
  assign statesOut_2_clock = clock;
  assign statesOut_2_reset = reset;
  assign statesOut_3_io_input_enable = swap;
  assign statesOut_3_clock = clock;
  assign statesOut_3_reset = reset;
  assign _T_164_data = io_input_0_data;
  assign _T_164_enable = _T_165;
  assign _T_164_reset = io_input_0_reset;
  assign _T_170_data = io_input_0_data;
  assign _T_170_enable = _T_171;
  assign _T_170_reset = io_input_0_reset;
  assign _T_176_data = io_input_0_data;
  assign _T_176_enable = _T_177;
  assign _T_176_reset = io_input_0_reset;
  assign _T_182_data = io_input_0_data;
  assign _T_182_enable = _T_183;
  assign _T_182_reset = io_input_0_reset;
  assign _T_226_0 = ff_0_io_output_data;
  assign _T_226_1 = ff_1_io_output_data;
  assign _T_226_2 = ff_2_io_output_data;
  assign _T_226_3 = ff_3_io_output_data;
  assign _T_246 = _T_244;
  assign _T_257_0 = ff_0_io_output_data;
  assign _T_257_1 = ff_1_io_output_data;
  assign _T_257_2 = ff_2_io_output_data;
  assign _T_257_3 = ff_3_io_output_data;
  assign _T_277 = _T_275;
  assign _T_288_0 = ff_0_io_output_data;
  assign _T_288_1 = ff_1_io_output_data;
  assign _T_288_2 = ff_2_io_output_data;
  assign _T_288_3 = ff_3_io_output_data;
  assign _T_308 = _T_306;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_149 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_149 <= 1'h0;
    end else begin
      _T_149 <= _T_146;
    end
  end
endmodule
module Mem1D(
  input         clock,
  input  [3:0]  io_w_addr,
  input  [31:0] io_w_data,
  input         io_w_en,
  input  [3:0]  io_r_addr,
  output [31:0] io_output_data
);
  reg [31:0] _T_14 [0:15];
  reg [31:0] _RAND_0;
  wire [31:0] _T_14__T_17_data;
  wire [3:0] _T_14__T_17_addr;
  wire [31:0] _T_14__T_16_data;
  wire [3:0] _T_14__T_16_addr;
  wire  _T_14__T_16_mask;
  wire  _T_14__T_16_en;
  assign _T_14__T_17_addr = io_r_addr;
  assign _T_14__T_17_data = _T_14[_T_14__T_17_addr];
  assign _T_14__T_16_data = io_w_data;
  assign _T_14__T_16_addr = io_w_addr;
  assign _T_14__T_16_mask = io_w_en;
  assign _T_14__T_16_en = io_w_en;
  assign io_output_data = _T_14__T_17_data;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    _T_14[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(_T_14__T_16_en & _T_14__T_16_mask) begin
      _T_14[_T_14__T_16_addr] <= _T_14__T_16_data;
    end
  end
endmodule
module MemND(
  input         clock,
  input  [3:0]  io_w_addr_0,
  input  [31:0] io_w_data,
  input         io_w_en,
  input         io_wMask,
  input  [3:0]  io_r_addr_0,
  output [31:0] io_output_data
);
  wire  m_clock;
  wire [3:0] m_io_w_addr;
  wire [31:0] m_io_w_data;
  wire  m_io_w_en;
  wire [3:0] m_io_r_addr;
  wire [31:0] m_io_output_data;
  wire [4:0] _T_17;
  wire [4:0] _T_20;
  wire  _T_22;
  Mem1D m (
    .clock(m_clock),
    .io_w_addr(m_io_w_addr),
    .io_w_data(m_io_w_data),
    .io_w_en(m_io_w_en),
    .io_r_addr(m_io_r_addr),
    .io_output_data(m_io_output_data)
  );
  assign _T_17 = io_w_addr_0 * 4'h1;
  assign _T_20 = io_r_addr_0 * 4'h1;
  assign _T_22 = io_w_en & io_wMask;
  assign io_output_data = m_io_output_data;
  assign m_io_w_addr = _T_17[3:0];
  assign m_io_w_data = io_w_data;
  assign m_io_w_en = _T_22;
  assign m_io_r_addr = _T_20[3:0];
  assign m_clock = clock;
endmodule
module SRAM(
  input         clock,
  input  [5:0]  io_w_0_addr_0,
  input  [31:0] io_w_0_data,
  input         io_w_0_en,
  input  [5:0]  io_r_0_addr_0,
  input         io_r_0_en,
  input  [5:0]  io_r_1_addr_0,
  input         io_r_1_en,
  input  [5:0]  io_r_2_addr_0,
  input         io_r_2_en,
  input  [5:0]  io_r_3_addr_0,
  output [31:0] io_output_data_0,
  output [31:0] io_output_data_1,
  output [31:0] io_output_data_2,
  output [31:0] io_output_data_3
);
  wire  m_0_clock;
  wire [3:0] m_0_io_w_addr_0;
  wire [31:0] m_0_io_w_data;
  wire  m_0_io_w_en;
  wire  m_0_io_wMask;
  wire [3:0] m_0_io_r_addr_0;
  wire [31:0] m_0_io_output_data;
  wire  m_1_clock;
  wire [3:0] m_1_io_w_addr_0;
  wire [31:0] m_1_io_w_data;
  wire  m_1_io_w_en;
  wire  m_1_io_wMask;
  wire [3:0] m_1_io_r_addr_0;
  wire [31:0] m_1_io_output_data;
  wire  m_2_clock;
  wire [3:0] m_2_io_w_addr_0;
  wire [31:0] m_2_io_w_data;
  wire  m_2_io_w_en;
  wire  m_2_io_wMask;
  wire [3:0] m_2_io_r_addr_0;
  wire [31:0] m_2_io_output_data;
  wire  m_3_clock;
  wire [3:0] m_3_io_w_addr_0;
  wire [31:0] m_3_io_w_data;
  wire  m_3_io_w_en;
  wire  m_3_io_wMask;
  wire [3:0] m_3_io_r_addr_0;
  wire [31:0] m_3_io_output_data;
  wire [5:0] convertedWVec_0_addr_0;
  wire [31:0] convertedWVec_0_data;
  wire  convertedWVec_0_en;
  wire [5:0] _T_35;
  wire [5:0] _GEN_0;
  wire [2:0] _T_37;
  wire [3:0] bankIdW_0;
  wire [5:0] convertedRVec_0_addr_0;
  wire  convertedRVec_0_en;
  wire [5:0] _T_43;
  wire [5:0] _GEN_1;
  wire [2:0] _T_46;
  wire [3:0] bankIdR_0;
  wire [5:0] convertedRVec_1_addr_0;
  wire  convertedRVec_1_en;
  wire [5:0] _T_52;
  wire [5:0] _GEN_2;
  wire [2:0] _T_55;
  wire [3:0] bankIdR_1;
  wire [5:0] convertedRVec_2_addr_0;
  wire  convertedRVec_2_en;
  wire [5:0] _T_61;
  wire [5:0] _GEN_3;
  wire [2:0] _T_64;
  wire [3:0] bankIdR_2;
  wire [5:0] convertedRVec_3_addr_0;
  wire [5:0] _T_70;
  wire [5:0] _GEN_4;
  wire [2:0] _T_73;
  wire [3:0] bankIdR_3;
  wire  _T_76;
  wire  _T_77;
  wire  _T_79;
  wire  _T_80;
  wire  _T_82;
  wire  _T_83;
  wire  _T_85;
  wire  _T_86;
  wire  _T_88;
  wire  _T_89;
  wire  _T_91;
  wire  _T_92;
  wire  _T_94;
  wire  _T_95;
  wire  _T_97;
  wire [5:0] _T_102_addr_0;
  wire [5:0] _T_104_addr_0;
  wire [5:0] _T_106_addr_0;
  wire  _T_109;
  wire  _T_110;
  wire  _T_112;
  wire  _T_113;
  wire  _T_115;
  wire  _T_116;
  wire  _T_118;
  wire [5:0] _T_123_addr_0;
  wire [5:0] _T_125_addr_0;
  wire [5:0] _T_127_addr_0;
  wire  _T_130;
  wire  _T_131;
  wire  _T_133;
  wire  _T_134;
  wire  _T_136;
  wire  _T_137;
  wire  _T_139;
  wire [5:0] _T_144_addr_0;
  wire [5:0] _T_146_addr_0;
  wire [5:0] _T_148_addr_0;
  wire  _T_151;
  wire  _T_152;
  wire  _T_154;
  wire  _T_155;
  wire  _T_157;
  wire  _T_158;
  wire [5:0] _T_165_addr_0;
  wire [5:0] _T_167_addr_0;
  wire [5:0] _T_169_addr_0;
  wire [31:0] _T_183;
  wire [31:0] _T_184;
  wire [31:0] _T_185;
  wire [31:0] _T_198;
  wire [31:0] _T_199;
  wire [31:0] _T_200;
  wire [31:0] _T_213;
  wire [31:0] _T_214;
  wire [31:0] _T_215;
  wire [31:0] _T_228;
  wire [31:0] _T_229;
  wire [31:0] _T_230;
  MemND m_0 (
    .clock(m_0_clock),
    .io_w_addr_0(m_0_io_w_addr_0),
    .io_w_data(m_0_io_w_data),
    .io_w_en(m_0_io_w_en),
    .io_wMask(m_0_io_wMask),
    .io_r_addr_0(m_0_io_r_addr_0),
    .io_output_data(m_0_io_output_data)
  );
  MemND m_1 (
    .clock(m_1_clock),
    .io_w_addr_0(m_1_io_w_addr_0),
    .io_w_data(m_1_io_w_data),
    .io_w_en(m_1_io_w_en),
    .io_wMask(m_1_io_wMask),
    .io_r_addr_0(m_1_io_r_addr_0),
    .io_output_data(m_1_io_output_data)
  );
  MemND m_2 (
    .clock(m_2_clock),
    .io_w_addr_0(m_2_io_w_addr_0),
    .io_w_data(m_2_io_w_data),
    .io_w_en(m_2_io_w_en),
    .io_wMask(m_2_io_wMask),
    .io_r_addr_0(m_2_io_r_addr_0),
    .io_output_data(m_2_io_output_data)
  );
  MemND m_3 (
    .clock(m_3_clock),
    .io_w_addr_0(m_3_io_w_addr_0),
    .io_w_data(m_3_io_w_data),
    .io_w_en(m_3_io_w_en),
    .io_wMask(m_3_io_wMask),
    .io_r_addr_0(m_3_io_r_addr_0),
    .io_output_data(m_3_io_output_data)
  );
  assign _T_35 = io_w_0_addr_0 / 6'h4;
  assign _GEN_0 = io_w_0_addr_0 % 6'h4;
  assign _T_37 = _GEN_0[2:0];
  assign bankIdW_0 = _T_37 * 3'h1;
  assign _T_43 = io_r_0_addr_0 / 6'h4;
  assign _GEN_1 = io_r_0_addr_0 % 6'h4;
  assign _T_46 = _GEN_1[2:0];
  assign bankIdR_0 = _T_46 * 3'h1;
  assign _T_52 = io_r_1_addr_0 / 6'h4;
  assign _GEN_2 = io_r_1_addr_0 % 6'h4;
  assign _T_55 = _GEN_2[2:0];
  assign bankIdR_1 = _T_55 * 3'h1;
  assign _T_61 = io_r_2_addr_0 / 6'h4;
  assign _GEN_3 = io_r_2_addr_0 % 6'h4;
  assign _T_64 = _GEN_3[2:0];
  assign bankIdR_2 = _T_64 * 3'h1;
  assign _T_70 = io_r_3_addr_0 / 6'h4;
  assign _GEN_4 = io_r_3_addr_0 % 6'h4;
  assign _T_73 = _GEN_4[2:0];
  assign bankIdR_3 = _T_73 * 3'h1;
  assign _T_76 = bankIdW_0 == 4'h0;
  assign _T_77 = _T_76 & convertedWVec_0_en;
  assign _T_79 = bankIdW_0 == 4'h1;
  assign _T_80 = _T_79 & convertedWVec_0_en;
  assign _T_82 = bankIdW_0 == 4'h2;
  assign _T_83 = _T_82 & convertedWVec_0_en;
  assign _T_85 = bankIdW_0 == 4'h3;
  assign _T_86 = _T_85 & convertedWVec_0_en;
  assign _T_88 = bankIdR_0 == 4'h0;
  assign _T_89 = _T_88 & convertedRVec_0_en;
  assign _T_91 = bankIdR_1 == 4'h0;
  assign _T_92 = _T_91 & convertedRVec_1_en;
  assign _T_94 = bankIdR_2 == 4'h0;
  assign _T_95 = _T_94 & convertedRVec_2_en;
  assign _T_97 = bankIdR_3 == 4'h0;
  assign _T_102_addr_0 = _T_95 ? convertedRVec_2_addr_0 : convertedRVec_3_addr_0;
  assign _T_104_addr_0 = _T_92 ? convertedRVec_1_addr_0 : _T_102_addr_0;
  assign _T_106_addr_0 = _T_89 ? convertedRVec_0_addr_0 : _T_104_addr_0;
  assign _T_109 = bankIdR_0 == 4'h1;
  assign _T_110 = _T_109 & convertedRVec_0_en;
  assign _T_112 = bankIdR_1 == 4'h1;
  assign _T_113 = _T_112 & convertedRVec_1_en;
  assign _T_115 = bankIdR_2 == 4'h1;
  assign _T_116 = _T_115 & convertedRVec_2_en;
  assign _T_118 = bankIdR_3 == 4'h1;
  assign _T_123_addr_0 = _T_116 ? convertedRVec_2_addr_0 : convertedRVec_3_addr_0;
  assign _T_125_addr_0 = _T_113 ? convertedRVec_1_addr_0 : _T_123_addr_0;
  assign _T_127_addr_0 = _T_110 ? convertedRVec_0_addr_0 : _T_125_addr_0;
  assign _T_130 = bankIdR_0 == 4'h2;
  assign _T_131 = _T_130 & convertedRVec_0_en;
  assign _T_133 = bankIdR_1 == 4'h2;
  assign _T_134 = _T_133 & convertedRVec_1_en;
  assign _T_136 = bankIdR_2 == 4'h2;
  assign _T_137 = _T_136 & convertedRVec_2_en;
  assign _T_139 = bankIdR_3 == 4'h2;
  assign _T_144_addr_0 = _T_137 ? convertedRVec_2_addr_0 : convertedRVec_3_addr_0;
  assign _T_146_addr_0 = _T_134 ? convertedRVec_1_addr_0 : _T_144_addr_0;
  assign _T_148_addr_0 = _T_131 ? convertedRVec_0_addr_0 : _T_146_addr_0;
  assign _T_151 = bankIdR_0 == 4'h3;
  assign _T_152 = _T_151 & convertedRVec_0_en;
  assign _T_154 = bankIdR_1 == 4'h3;
  assign _T_155 = _T_154 & convertedRVec_1_en;
  assign _T_157 = bankIdR_2 == 4'h3;
  assign _T_158 = _T_157 & convertedRVec_2_en;
  assign _T_165_addr_0 = _T_158 ? convertedRVec_2_addr_0 : convertedRVec_3_addr_0;
  assign _T_167_addr_0 = _T_155 ? convertedRVec_1_addr_0 : _T_165_addr_0;
  assign _T_169_addr_0 = _T_152 ? convertedRVec_0_addr_0 : _T_167_addr_0;
  assign _T_183 = _T_130 ? m_2_io_output_data : m_3_io_output_data;
  assign _T_184 = _T_109 ? m_1_io_output_data : _T_183;
  assign _T_185 = _T_88 ? m_0_io_output_data : _T_184;
  assign _T_198 = _T_133 ? m_2_io_output_data : m_3_io_output_data;
  assign _T_199 = _T_112 ? m_1_io_output_data : _T_198;
  assign _T_200 = _T_91 ? m_0_io_output_data : _T_199;
  assign _T_213 = _T_136 ? m_2_io_output_data : m_3_io_output_data;
  assign _T_214 = _T_115 ? m_1_io_output_data : _T_213;
  assign _T_215 = _T_94 ? m_0_io_output_data : _T_214;
  assign _T_228 = _T_139 ? m_2_io_output_data : m_3_io_output_data;
  assign _T_229 = _T_118 ? m_1_io_output_data : _T_228;
  assign _T_230 = _T_97 ? m_0_io_output_data : _T_229;
  assign io_output_data_0 = _T_185;
  assign io_output_data_1 = _T_200;
  assign io_output_data_2 = _T_215;
  assign io_output_data_3 = _T_230;
  assign m_0_io_w_addr_0 = convertedWVec_0_addr_0[3:0];
  assign m_0_io_w_data = convertedWVec_0_data;
  assign m_0_io_w_en = convertedWVec_0_en;
  assign m_0_io_wMask = _T_77;
  assign m_0_io_r_addr_0 = _T_106_addr_0[3:0];
  assign m_0_clock = clock;
  assign m_1_io_w_addr_0 = convertedWVec_0_addr_0[3:0];
  assign m_1_io_w_data = convertedWVec_0_data;
  assign m_1_io_w_en = convertedWVec_0_en;
  assign m_1_io_wMask = _T_80;
  assign m_1_io_r_addr_0 = _T_127_addr_0[3:0];
  assign m_1_clock = clock;
  assign m_2_io_w_addr_0 = convertedWVec_0_addr_0[3:0];
  assign m_2_io_w_data = convertedWVec_0_data;
  assign m_2_io_w_en = convertedWVec_0_en;
  assign m_2_io_wMask = _T_83;
  assign m_2_io_r_addr_0 = _T_148_addr_0[3:0];
  assign m_2_clock = clock;
  assign m_3_io_w_addr_0 = convertedWVec_0_addr_0[3:0];
  assign m_3_io_w_data = convertedWVec_0_data;
  assign m_3_io_w_en = convertedWVec_0_en;
  assign m_3_io_wMask = _T_86;
  assign m_3_io_r_addr_0 = _T_169_addr_0[3:0];
  assign m_3_clock = clock;
  assign convertedWVec_0_addr_0 = _T_35;
  assign convertedWVec_0_data = io_w_0_data;
  assign convertedWVec_0_en = io_w_0_en;
  assign convertedRVec_0_addr_0 = _T_43;
  assign convertedRVec_0_en = io_r_0_en;
  assign convertedRVec_1_addr_0 = _T_52;
  assign convertedRVec_1_en = io_r_1_en;
  assign convertedRVec_2_addr_0 = _T_61;
  assign convertedRVec_2_en = io_r_2_en;
  assign convertedRVec_3_addr_0 = _T_70;
endmodule
module NBufCtr_22(
  input        clock,
  input        reset,
  input        io_input_countUp,
  input        io_input_enable,
  output [2:0] io_output_count
);
  wire [2:0] _T_8;
  wire [3:0] _T_10;
  wire [2:0] _T_11;
  wire  _T_13;
  wire [2:0] _T_14;
  wire [3:0] _T_16;
  wire [2:0] _T_17;
  wire [2:0] _T_18;
  wire [2:0] _T_19;
  wire [2:0] _T_23;
  wire  _T_25;
  wire [3:0] _T_28;
  wire [3:0] _T_29;
  wire [2:0] _T_30;
  wire [2:0] _T_31;
  wire [2:0] _T_32;
  wire [3:0] _T_34;
  wire [2:0] _T_35;
  wire  _T_37;
  wire [3:0] _T_41;
  wire [2:0] _T_42;
  wire [2:0] _T_43;
  wire [2:0] _T_44;
  wire [3:0] _T_45;
  wire [2:0] _T_46;
  wire [2:0] _T_50;
  wire [2:0] _T_51;
  wire [2:0] _T_54;
  wire [2:0] _T_55;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire [2:0] RetimeWrapper_io_in;
  wire [2:0] RetimeWrapper_io_out;
  wire [2:0] _T_59;
  RetimeWrapper_106 RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_10 = _T_8 + 3'h0;
  assign _T_11 = _T_10[2:0];
  assign _T_13 = _T_11 >= 3'h3;
  assign _T_14 = $signed(_T_8);
  assign _T_16 = $signed(_T_14) + $signed(-3'sh3);
  assign _T_17 = _T_16[2:0];
  assign _T_18 = $signed(_T_17);
  assign _T_19 = $unsigned(_T_18);
  assign _T_23 = _T_13 ? _T_19 : _T_11;
  assign _T_25 = _T_8 == 3'h0;
  assign _T_28 = _T_8 - 3'h1;
  assign _T_29 = $unsigned(_T_28);
  assign _T_30 = _T_29[2:0];
  assign _T_31 = _T_25 ? 3'h2 : _T_30;
  assign _T_32 = io_input_enable ? _T_31 : _T_8;
  assign _T_34 = _T_8 + 3'h1;
  assign _T_35 = _T_34[2:0];
  assign _T_37 = _T_35 >= 3'h3;
  assign _T_41 = $signed(_T_14) + $signed(-3'sh2);
  assign _T_42 = _T_41[2:0];
  assign _T_43 = $signed(_T_42);
  assign _T_44 = $unsigned(_T_43);
  assign _T_45 = 3'h0 + _T_44;
  assign _T_46 = _T_45[2:0];
  assign _T_50 = _T_37 ? _T_46 : _T_35;
  assign _T_51 = io_input_enable ? _T_50 : _T_8;
  assign _T_54 = io_input_countUp ? _T_51 : _T_32;
  assign _T_55 = reset ? 3'h0 : _T_54;
  assign io_output_count = _T_23;
  assign _T_8 = _T_59;
  assign RetimeWrapper_io_in = _T_55;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_59 = RetimeWrapper_io_out;
endmodule
module NBufCtr_24(
  input        clock,
  input        reset,
  input        io_input_countUp,
  input        io_input_enable,
  output [2:0] io_output_count
);
  wire [2:0] _T_8;
  wire [3:0] _T_10;
  wire [2:0] _T_11;
  wire  _T_13;
  wire [2:0] _T_14;
  wire [3:0] _T_16;
  wire [2:0] _T_17;
  wire [2:0] _T_18;
  wire [2:0] _T_19;
  wire [2:0] _T_23;
  wire  _T_25;
  wire [3:0] _T_28;
  wire [3:0] _T_29;
  wire [2:0] _T_30;
  wire [2:0] _T_31;
  wire [2:0] _T_32;
  wire [3:0] _T_45;
  wire [2:0] _T_46;
  wire [2:0] _T_50;
  wire [2:0] _T_51;
  wire [2:0] _T_54;
  wire [2:0] _T_55;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire [2:0] RetimeWrapper_io_in;
  wire [2:0] RetimeWrapper_io_out;
  wire [2:0] _T_59;
  RetimeWrapper_106 RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_10 = _T_8 + 3'h1;
  assign _T_11 = _T_10[2:0];
  assign _T_13 = _T_11 >= 3'h3;
  assign _T_14 = $signed(_T_8);
  assign _T_16 = $signed(_T_14) + $signed(-3'sh2);
  assign _T_17 = _T_16[2:0];
  assign _T_18 = $signed(_T_17);
  assign _T_19 = $unsigned(_T_18);
  assign _T_23 = _T_13 ? _T_19 : _T_11;
  assign _T_25 = _T_8 == 3'h0;
  assign _T_28 = _T_8 - 3'h1;
  assign _T_29 = $unsigned(_T_28);
  assign _T_30 = _T_29[2:0];
  assign _T_31 = _T_25 ? 3'h2 : _T_30;
  assign _T_32 = io_input_enable ? _T_31 : _T_8;
  assign _T_45 = 3'h0 + _T_19;
  assign _T_46 = _T_45[2:0];
  assign _T_50 = _T_13 ? _T_46 : _T_11;
  assign _T_51 = io_input_enable ? _T_50 : _T_8;
  assign _T_54 = io_input_countUp ? _T_51 : _T_32;
  assign _T_55 = reset ? 3'h0 : _T_54;
  assign io_output_count = _T_23;
  assign _T_8 = _T_59;
  assign RetimeWrapper_io_in = _T_55;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_59 = RetimeWrapper_io_out;
endmodule
module NBufCtr_25(
  input        clock,
  input        reset,
  input        io_input_countUp,
  input        io_input_enable,
  output [2:0] io_output_count
);
  wire [2:0] _T_8;
  wire [3:0] _T_10;
  wire [2:0] _T_11;
  wire  _T_13;
  wire [2:0] _T_14;
  wire [3:0] _T_16;
  wire [2:0] _T_17;
  wire [2:0] _T_18;
  wire [2:0] _T_19;
  wire [2:0] _T_23;
  wire  _T_25;
  wire [3:0] _T_28;
  wire [3:0] _T_29;
  wire [2:0] _T_30;
  wire [2:0] _T_31;
  wire [2:0] _T_32;
  wire [3:0] _T_34;
  wire [2:0] _T_35;
  wire  _T_37;
  wire [3:0] _T_41;
  wire [2:0] _T_42;
  wire [2:0] _T_43;
  wire [2:0] _T_44;
  wire [3:0] _T_45;
  wire [2:0] _T_46;
  wire [2:0] _T_50;
  wire [2:0] _T_51;
  wire [2:0] _T_54;
  wire [2:0] _T_55;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire [2:0] RetimeWrapper_io_in;
  wire [2:0] RetimeWrapper_io_out;
  wire [2:0] _T_59;
  RetimeWrapper_106 RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_10 = _T_8 + 3'h2;
  assign _T_11 = _T_10[2:0];
  assign _T_13 = _T_11 >= 3'h3;
  assign _T_14 = $signed(_T_8);
  assign _T_16 = $signed(_T_14) + $signed(-3'sh1);
  assign _T_17 = _T_16[2:0];
  assign _T_18 = $signed(_T_17);
  assign _T_19 = $unsigned(_T_18);
  assign _T_23 = _T_13 ? _T_19 : _T_11;
  assign _T_25 = _T_8 == 3'h0;
  assign _T_28 = _T_8 - 3'h1;
  assign _T_29 = $unsigned(_T_28);
  assign _T_30 = _T_29[2:0];
  assign _T_31 = _T_25 ? 3'h2 : _T_30;
  assign _T_32 = io_input_enable ? _T_31 : _T_8;
  assign _T_34 = _T_8 + 3'h1;
  assign _T_35 = _T_34[2:0];
  assign _T_37 = _T_35 >= 3'h3;
  assign _T_41 = $signed(_T_14) + $signed(-3'sh2);
  assign _T_42 = _T_41[2:0];
  assign _T_43 = $signed(_T_42);
  assign _T_44 = $unsigned(_T_43);
  assign _T_45 = 3'h0 + _T_44;
  assign _T_46 = _T_45[2:0];
  assign _T_50 = _T_37 ? _T_46 : _T_35;
  assign _T_51 = io_input_enable ? _T_50 : _T_8;
  assign _T_54 = io_input_countUp ? _T_51 : _T_32;
  assign _T_55 = reset ? 3'h0 : _T_54;
  assign io_output_count = _T_23;
  assign _T_8 = _T_59;
  assign RetimeWrapper_io_in = _T_55;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_59 = RetimeWrapper_io_out;
endmodule
module NBufSRAMnoBcast(
  input         clock,
  input         reset,
  input         io_sEn_0,
  input         io_sEn_1,
  input         io_sEn_2,
  input         io_sDone_0,
  input         io_sDone_1,
  input         io_sDone_2,
  input  [5:0]  io_w_0_addr_0,
  input  [31:0] io_w_0_data,
  input         io_w_0_en,
  input  [5:0]  io_r_0_addr_0,
  input         io_r_0_en,
  input  [5:0]  io_r_1_addr_0,
  input         io_r_1_en,
  input  [5:0]  io_r_2_addr_0,
  input         io_r_2_en,
  input  [5:0]  io_r_3_addr_0,
  input         io_r_3_en,
  output [31:0] io_output_data_8,
  output [31:0] io_output_data_9,
  output [31:0] io_output_data_10,
  output [31:0] io_output_data_11
);
  wire  srams_0_clock;
  wire [5:0] srams_0_io_w_0_addr_0;
  wire [31:0] srams_0_io_w_0_data;
  wire  srams_0_io_w_0_en;
  wire [5:0] srams_0_io_r_0_addr_0;
  wire  srams_0_io_r_0_en;
  wire [5:0] srams_0_io_r_1_addr_0;
  wire  srams_0_io_r_1_en;
  wire [5:0] srams_0_io_r_2_addr_0;
  wire  srams_0_io_r_2_en;
  wire [5:0] srams_0_io_r_3_addr_0;
  wire [31:0] srams_0_io_output_data_0;
  wire [31:0] srams_0_io_output_data_1;
  wire [31:0] srams_0_io_output_data_2;
  wire [31:0] srams_0_io_output_data_3;
  wire  srams_1_clock;
  wire [5:0] srams_1_io_w_0_addr_0;
  wire [31:0] srams_1_io_w_0_data;
  wire  srams_1_io_w_0_en;
  wire [5:0] srams_1_io_r_0_addr_0;
  wire  srams_1_io_r_0_en;
  wire [5:0] srams_1_io_r_1_addr_0;
  wire  srams_1_io_r_1_en;
  wire [5:0] srams_1_io_r_2_addr_0;
  wire  srams_1_io_r_2_en;
  wire [5:0] srams_1_io_r_3_addr_0;
  wire [31:0] srams_1_io_output_data_0;
  wire [31:0] srams_1_io_output_data_1;
  wire [31:0] srams_1_io_output_data_2;
  wire [31:0] srams_1_io_output_data_3;
  wire  srams_2_clock;
  wire [5:0] srams_2_io_w_0_addr_0;
  wire [31:0] srams_2_io_w_0_data;
  wire  srams_2_io_w_0_en;
  wire [5:0] srams_2_io_r_0_addr_0;
  wire  srams_2_io_r_0_en;
  wire [5:0] srams_2_io_r_1_addr_0;
  wire  srams_2_io_r_1_en;
  wire [5:0] srams_2_io_r_2_addr_0;
  wire  srams_2_io_r_2_en;
  wire [5:0] srams_2_io_r_3_addr_0;
  wire [31:0] srams_2_io_output_data_0;
  wire [31:0] srams_2_io_output_data_1;
  wire [31:0] srams_2_io_output_data_2;
  wire [31:0] srams_2_io_output_data_3;
  wire  sEn_latch_0_clock;
  wire  sEn_latch_0_reset;
  wire  sEn_latch_0_io_input_set;
  wire  sEn_latch_0_io_input_reset;
  wire  sEn_latch_0_io_input_asyn_reset;
  wire  sEn_latch_0_io_output_data;
  wire  sEn_latch_1_clock;
  wire  sEn_latch_1_reset;
  wire  sEn_latch_1_io_input_set;
  wire  sEn_latch_1_io_input_reset;
  wire  sEn_latch_1_io_input_asyn_reset;
  wire  sEn_latch_1_io_output_data;
  wire  sEn_latch_2_clock;
  wire  sEn_latch_2_reset;
  wire  sEn_latch_2_io_input_set;
  wire  sEn_latch_2_io_input_reset;
  wire  sEn_latch_2_io_input_asyn_reset;
  wire  sEn_latch_2_io_output_data;
  wire  sDone_latch_0_clock;
  wire  sDone_latch_0_reset;
  wire  sDone_latch_0_io_input_set;
  wire  sDone_latch_0_io_input_reset;
  wire  sDone_latch_0_io_input_asyn_reset;
  wire  sDone_latch_0_io_output_data;
  wire  sDone_latch_1_clock;
  wire  sDone_latch_1_reset;
  wire  sDone_latch_1_io_input_set;
  wire  sDone_latch_1_io_input_reset;
  wire  sDone_latch_1_io_input_asyn_reset;
  wire  sDone_latch_1_io_output_data;
  wire  sDone_latch_2_clock;
  wire  sDone_latch_2_reset;
  wire  sDone_latch_2_io_input_set;
  wire  sDone_latch_2_io_input_reset;
  wire  sDone_latch_2_io_input_asyn_reset;
  wire  sDone_latch_2_io_output_data;
  wire  swap;
  wire  _T_38;
  wire  _T_39;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire  RetimeWrapper_io_flow;
  wire  RetimeWrapper_io_in;
  wire  RetimeWrapper_io_out;
  wire  _T_43;
  wire  RetimeWrapper_1_clock;
  wire  RetimeWrapper_1_reset;
  wire  RetimeWrapper_1_io_flow;
  wire  RetimeWrapper_1_io_in;
  wire  RetimeWrapper_1_io_out;
  wire  _T_47;
  wire  RetimeWrapper_2_clock;
  wire  RetimeWrapper_2_reset;
  wire  RetimeWrapper_2_io_flow;
  wire  RetimeWrapper_2_io_in;
  wire  RetimeWrapper_2_io_out;
  wire  _T_51;
  wire  RetimeWrapper_3_clock;
  wire  RetimeWrapper_3_reset;
  wire  RetimeWrapper_3_io_flow;
  wire  RetimeWrapper_3_io_in;
  wire  RetimeWrapper_3_io_out;
  wire  _T_55;
  wire  _T_56;
  wire  _T_57;
  wire  RetimeWrapper_4_clock;
  wire  RetimeWrapper_4_reset;
  wire  RetimeWrapper_4_io_flow;
  wire  RetimeWrapper_4_io_in;
  wire  RetimeWrapper_4_io_out;
  wire  _T_61;
  wire  RetimeWrapper_5_clock;
  wire  RetimeWrapper_5_reset;
  wire  RetimeWrapper_5_io_flow;
  wire  RetimeWrapper_5_io_in;
  wire  RetimeWrapper_5_io_out;
  wire  _T_65;
  wire  RetimeWrapper_6_clock;
  wire  RetimeWrapper_6_reset;
  wire  RetimeWrapper_6_io_flow;
  wire  RetimeWrapper_6_io_in;
  wire  RetimeWrapper_6_io_out;
  wire  _T_69;
  wire  RetimeWrapper_7_clock;
  wire  RetimeWrapper_7_reset;
  wire  RetimeWrapper_7_io_flow;
  wire  RetimeWrapper_7_io_in;
  wire  RetimeWrapper_7_io_out;
  wire  _T_73;
  wire  _T_74;
  wire  _T_75;
  wire  RetimeWrapper_8_clock;
  wire  RetimeWrapper_8_reset;
  wire  RetimeWrapper_8_io_flow;
  wire  RetimeWrapper_8_io_in;
  wire  RetimeWrapper_8_io_out;
  wire  _T_79;
  wire  RetimeWrapper_9_clock;
  wire  RetimeWrapper_9_reset;
  wire  RetimeWrapper_9_io_flow;
  wire  RetimeWrapper_9_io_in;
  wire  RetimeWrapper_9_io_out;
  wire  _T_83;
  wire  RetimeWrapper_10_clock;
  wire  RetimeWrapper_10_reset;
  wire  RetimeWrapper_10_io_flow;
  wire  RetimeWrapper_10_io_in;
  wire  RetimeWrapper_10_io_out;
  wire  _T_87;
  wire  RetimeWrapper_11_clock;
  wire  RetimeWrapper_11_reset;
  wire  RetimeWrapper_11_io_flow;
  wire  RetimeWrapper_11_io_in;
  wire  RetimeWrapper_11_io_out;
  wire  _T_91;
  wire  _T_92;
  wire  anyEnabled;
  wire  _T_93;
  wire  _T_94;
  wire  _T_95;
  wire  _T_96;
  wire  _T_97;
  wire  _T_98;
  wire  _T_99;
  wire  _T_100;
  wire  _T_101;
  wire  _T_102;
  reg  _T_105;
  reg [31:0] _RAND_0;
  wire  _T_111;
  wire  NBufCtr_clock;
  wire  NBufCtr_reset;
  wire  NBufCtr_io_input_countUp;
  wire  NBufCtr_io_input_enable;
  wire [2:0] NBufCtr_io_output_count;
  wire  statesInR_0_clock;
  wire  statesInR_0_reset;
  wire  statesInR_0_io_input_countUp;
  wire  statesInR_0_io_input_enable;
  wire [2:0] statesInR_0_io_output_count;
  wire  statesInR_1_clock;
  wire  statesInR_1_reset;
  wire  statesInR_1_io_input_countUp;
  wire  statesInR_1_io_input_enable;
  wire [2:0] statesInR_1_io_output_count;
  wire  statesInR_2_clock;
  wire  statesInR_2_reset;
  wire  statesInR_2_io_input_countUp;
  wire  statesInR_2_io_input_enable;
  wire [2:0] statesInR_2_io_output_count;
  wire  statesOut_0_clock;
  wire  statesOut_0_reset;
  wire  statesOut_0_io_input_countUp;
  wire  statesOut_0_io_input_enable;
  wire [2:0] statesOut_0_io_output_count;
  wire  statesOut_1_clock;
  wire  statesOut_1_reset;
  wire  statesOut_1_io_input_countUp;
  wire  statesOut_1_io_input_enable;
  wire [2:0] statesOut_1_io_output_count;
  wire  statesOut_2_clock;
  wire  statesOut_2_reset;
  wire  statesOut_2_io_input_countUp;
  wire  statesOut_2_io_input_enable;
  wire [2:0] statesOut_2_io_output_count;
  wire  _T_120;
  wire [5:0] _T_124_addr_0;
  wire [31:0] _T_124_data;
  wire  _T_124_en;
  wire  _T_126;
  wire  _T_134;
  wire [6:0] _T_159;
  wire [6:0] _T_161;
  wire [5:0] _T_166_addr_0;
  wire  _T_166_en;
  wire [6:0] _T_169;
  wire  _T_170;
  wire [5:0] _T_171;
  wire [6:0] _T_195;
  wire [6:0] _T_197;
  wire [5:0] _T_202_addr_0;
  wire  _T_202_en;
  wire [6:0] _T_205;
  wire  _T_206;
  wire [5:0] _T_207;
  wire [6:0] _T_231;
  wire [6:0] _T_233;
  wire [5:0] _T_238_addr_0;
  wire  _T_238_en;
  wire [6:0] _T_241;
  wire  _T_242;
  wire [5:0] _T_243;
  wire [6:0] _T_267;
  wire [6:0] _T_269;
  wire [5:0] _T_274_addr_0;
  wire [6:0] _T_277;
  wire [5:0] _T_279;
  wire  _T_281;
  wire [5:0] _T_285_addr_0;
  wire [31:0] _T_285_data;
  wire  _T_285_en;
  wire  _T_287;
  wire  _T_295;
  wire [6:0] _T_322;
  wire [5:0] _T_327_addr_0;
  wire  _T_327_en;
  wire [6:0] _T_330;
  wire  _T_331;
  wire [5:0] _T_332;
  wire [6:0] _T_358;
  wire [5:0] _T_363_addr_0;
  wire  _T_363_en;
  wire [6:0] _T_366;
  wire  _T_367;
  wire [5:0] _T_368;
  wire [6:0] _T_394;
  wire [5:0] _T_399_addr_0;
  wire  _T_399_en;
  wire [6:0] _T_402;
  wire  _T_403;
  wire [5:0] _T_404;
  wire [6:0] _T_430;
  wire [5:0] _T_435_addr_0;
  wire [6:0] _T_438;
  wire [5:0] _T_440;
  wire  _T_442;
  wire [5:0] _T_446_addr_0;
  wire [31:0] _T_446_data;
  wire  _T_446_en;
  wire  _T_448;
  wire  _T_456;
  wire [6:0] _T_483;
  wire [5:0] _T_488_addr_0;
  wire  _T_488_en;
  wire [6:0] _T_491;
  wire  _T_492;
  wire [5:0] _T_493;
  wire [6:0] _T_519;
  wire [5:0] _T_524_addr_0;
  wire  _T_524_en;
  wire [6:0] _T_527;
  wire  _T_528;
  wire [5:0] _T_529;
  wire [6:0] _T_555;
  wire [5:0] _T_560_addr_0;
  wire  _T_560_en;
  wire [6:0] _T_563;
  wire  _T_564;
  wire [5:0] _T_565;
  wire [6:0] _T_591;
  wire [5:0] _T_596_addr_0;
  wire [6:0] _T_599;
  wire [5:0] _T_601;
  wire  _T_709;
  wire  _T_712;
  wire  _T_715;
  wire [31:0] _T_719;
  wire [31:0] _T_721;
  wire [31:0] _T_723;
  wire [31:0] _T_724;
  wire [31:0] _T_725;
  wire [31:0] _T_727;
  wire [31:0] _T_730;
  wire [31:0] _T_732;
  wire [31:0] _T_734;
  wire [31:0] _T_735;
  wire [31:0] _T_736;
  wire [31:0] _T_738;
  wire [31:0] _T_741;
  wire [31:0] _T_743;
  wire [31:0] _T_745;
  wire [31:0] _T_746;
  wire [31:0] _T_747;
  wire [31:0] _T_749;
  wire [31:0] _T_752;
  wire [31:0] _T_754;
  wire [31:0] _T_756;
  wire [31:0] _T_757;
  wire [31:0] _T_758;
  wire [31:0] _T_760;
  SRAM srams_0 (
    .clock(srams_0_clock),
    .io_w_0_addr_0(srams_0_io_w_0_addr_0),
    .io_w_0_data(srams_0_io_w_0_data),
    .io_w_0_en(srams_0_io_w_0_en),
    .io_r_0_addr_0(srams_0_io_r_0_addr_0),
    .io_r_0_en(srams_0_io_r_0_en),
    .io_r_1_addr_0(srams_0_io_r_1_addr_0),
    .io_r_1_en(srams_0_io_r_1_en),
    .io_r_2_addr_0(srams_0_io_r_2_addr_0),
    .io_r_2_en(srams_0_io_r_2_en),
    .io_r_3_addr_0(srams_0_io_r_3_addr_0),
    .io_output_data_0(srams_0_io_output_data_0),
    .io_output_data_1(srams_0_io_output_data_1),
    .io_output_data_2(srams_0_io_output_data_2),
    .io_output_data_3(srams_0_io_output_data_3)
  );
  SRAM srams_1 (
    .clock(srams_1_clock),
    .io_w_0_addr_0(srams_1_io_w_0_addr_0),
    .io_w_0_data(srams_1_io_w_0_data),
    .io_w_0_en(srams_1_io_w_0_en),
    .io_r_0_addr_0(srams_1_io_r_0_addr_0),
    .io_r_0_en(srams_1_io_r_0_en),
    .io_r_1_addr_0(srams_1_io_r_1_addr_0),
    .io_r_1_en(srams_1_io_r_1_en),
    .io_r_2_addr_0(srams_1_io_r_2_addr_0),
    .io_r_2_en(srams_1_io_r_2_en),
    .io_r_3_addr_0(srams_1_io_r_3_addr_0),
    .io_output_data_0(srams_1_io_output_data_0),
    .io_output_data_1(srams_1_io_output_data_1),
    .io_output_data_2(srams_1_io_output_data_2),
    .io_output_data_3(srams_1_io_output_data_3)
  );
  SRAM srams_2 (
    .clock(srams_2_clock),
    .io_w_0_addr_0(srams_2_io_w_0_addr_0),
    .io_w_0_data(srams_2_io_w_0_data),
    .io_w_0_en(srams_2_io_w_0_en),
    .io_r_0_addr_0(srams_2_io_r_0_addr_0),
    .io_r_0_en(srams_2_io_r_0_en),
    .io_r_1_addr_0(srams_2_io_r_1_addr_0),
    .io_r_1_en(srams_2_io_r_1_en),
    .io_r_2_addr_0(srams_2_io_r_2_addr_0),
    .io_r_2_en(srams_2_io_r_2_en),
    .io_r_3_addr_0(srams_2_io_r_3_addr_0),
    .io_output_data_0(srams_2_io_output_data_0),
    .io_output_data_1(srams_2_io_output_data_1),
    .io_output_data_2(srams_2_io_output_data_2),
    .io_output_data_3(srams_2_io_output_data_3)
  );
  SRFF sEn_latch_0 (
    .clock(sEn_latch_0_clock),
    .reset(sEn_latch_0_reset),
    .io_input_set(sEn_latch_0_io_input_set),
    .io_input_reset(sEn_latch_0_io_input_reset),
    .io_input_asyn_reset(sEn_latch_0_io_input_asyn_reset),
    .io_output_data(sEn_latch_0_io_output_data)
  );
  SRFF sEn_latch_1 (
    .clock(sEn_latch_1_clock),
    .reset(sEn_latch_1_reset),
    .io_input_set(sEn_latch_1_io_input_set),
    .io_input_reset(sEn_latch_1_io_input_reset),
    .io_input_asyn_reset(sEn_latch_1_io_input_asyn_reset),
    .io_output_data(sEn_latch_1_io_output_data)
  );
  SRFF sEn_latch_2 (
    .clock(sEn_latch_2_clock),
    .reset(sEn_latch_2_reset),
    .io_input_set(sEn_latch_2_io_input_set),
    .io_input_reset(sEn_latch_2_io_input_reset),
    .io_input_asyn_reset(sEn_latch_2_io_input_asyn_reset),
    .io_output_data(sEn_latch_2_io_output_data)
  );
  SRFF sDone_latch_0 (
    .clock(sDone_latch_0_clock),
    .reset(sDone_latch_0_reset),
    .io_input_set(sDone_latch_0_io_input_set),
    .io_input_reset(sDone_latch_0_io_input_reset),
    .io_input_asyn_reset(sDone_latch_0_io_input_asyn_reset),
    .io_output_data(sDone_latch_0_io_output_data)
  );
  SRFF sDone_latch_1 (
    .clock(sDone_latch_1_clock),
    .reset(sDone_latch_1_reset),
    .io_input_set(sDone_latch_1_io_input_set),
    .io_input_reset(sDone_latch_1_io_input_reset),
    .io_input_asyn_reset(sDone_latch_1_io_input_asyn_reset),
    .io_output_data(sDone_latch_1_io_output_data)
  );
  SRFF sDone_latch_2 (
    .clock(sDone_latch_2_clock),
    .reset(sDone_latch_2_reset),
    .io_input_set(sDone_latch_2_io_input_set),
    .io_input_reset(sDone_latch_2_io_input_reset),
    .io_input_asyn_reset(sDone_latch_2_io_input_asyn_reset),
    .io_output_data(sDone_latch_2_io_output_data)
  );
  RetimeWrapper RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 (
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 (
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 (
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 (
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 (
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 (
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 (
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper RetimeWrapper_8 (
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper RetimeWrapper_9 (
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper RetimeWrapper_10 (
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper RetimeWrapper_11 (
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  NBufCtr_22 NBufCtr (
    .clock(NBufCtr_clock),
    .reset(NBufCtr_reset),
    .io_input_countUp(NBufCtr_io_input_countUp),
    .io_input_enable(NBufCtr_io_input_enable),
    .io_output_count(NBufCtr_io_output_count)
  );
  NBufCtr_22 statesInR_0 (
    .clock(statesInR_0_clock),
    .reset(statesInR_0_reset),
    .io_input_countUp(statesInR_0_io_input_countUp),
    .io_input_enable(statesInR_0_io_input_enable),
    .io_output_count(statesInR_0_io_output_count)
  );
  NBufCtr_24 statesInR_1 (
    .clock(statesInR_1_clock),
    .reset(statesInR_1_reset),
    .io_input_countUp(statesInR_1_io_input_countUp),
    .io_input_enable(statesInR_1_io_input_enable),
    .io_output_count(statesInR_1_io_output_count)
  );
  NBufCtr_25 statesInR_2 (
    .clock(statesInR_2_clock),
    .reset(statesInR_2_reset),
    .io_input_countUp(statesInR_2_io_input_countUp),
    .io_input_enable(statesInR_2_io_input_enable),
    .io_output_count(statesInR_2_io_output_count)
  );
  NBufCtr_22 statesOut_0 (
    .clock(statesOut_0_clock),
    .reset(statesOut_0_reset),
    .io_input_countUp(statesOut_0_io_input_countUp),
    .io_input_enable(statesOut_0_io_input_enable),
    .io_output_count(statesOut_0_io_output_count)
  );
  NBufCtr_24 statesOut_1 (
    .clock(statesOut_1_clock),
    .reset(statesOut_1_reset),
    .io_input_countUp(statesOut_1_io_input_countUp),
    .io_input_enable(statesOut_1_io_input_enable),
    .io_output_count(statesOut_1_io_output_count)
  );
  NBufCtr_25 statesOut_2 (
    .clock(statesOut_2_clock),
    .reset(statesOut_2_reset),
    .io_input_countUp(statesOut_2_io_input_countUp),
    .io_input_enable(statesOut_2_io_input_enable),
    .io_output_count(statesOut_2_io_output_count)
  );
  assign _T_38 = ~ io_sDone_0;
  assign _T_39 = io_sEn_0 & _T_38;
  assign _T_56 = ~ io_sDone_1;
  assign _T_57 = io_sEn_1 & _T_56;
  assign _T_74 = ~ io_sDone_2;
  assign _T_75 = io_sEn_2 & _T_74;
  assign _T_92 = sEn_latch_0_io_output_data | sEn_latch_1_io_output_data;
  assign anyEnabled = _T_92 | sEn_latch_2_io_output_data;
  assign _T_93 = sDone_latch_0_io_output_data | io_sDone_0;
  assign _T_94 = sEn_latch_0_io_output_data == _T_93;
  assign _T_95 = sDone_latch_1_io_output_data | io_sDone_1;
  assign _T_96 = sEn_latch_1_io_output_data == _T_95;
  assign _T_97 = sDone_latch_2_io_output_data | io_sDone_2;
  assign _T_98 = sEn_latch_2_io_output_data == _T_97;
  assign _T_99 = _T_94 & _T_96;
  assign _T_100 = _T_99 & _T_98;
  assign _T_101 = _T_100 & anyEnabled;
  assign _T_102 = ~ _T_101;
  assign _T_111 = _T_101 & _T_105;
  assign _T_120 = NBufCtr_io_output_count == 3'h0;
  assign _T_126 = io_w_0_en & _T_120;
  assign _T_134 = statesInR_0_io_output_count == 3'h2;
  assign _T_159 = {io_r_0_addr_0,io_r_0_en};
  assign _T_161 = _T_134 ? _T_159 : 7'h0;
  assign _T_170 = _T_169[0];
  assign _T_171 = _T_169[6:1];
  assign _T_195 = {io_r_1_addr_0,io_r_1_en};
  assign _T_197 = _T_134 ? _T_195 : 7'h0;
  assign _T_206 = _T_205[0];
  assign _T_207 = _T_205[6:1];
  assign _T_231 = {io_r_2_addr_0,io_r_2_en};
  assign _T_233 = _T_134 ? _T_231 : 7'h0;
  assign _T_242 = _T_241[0];
  assign _T_243 = _T_241[6:1];
  assign _T_267 = {io_r_3_addr_0,io_r_3_en};
  assign _T_269 = _T_134 ? _T_267 : 7'h0;
  assign _T_279 = _T_277[6:1];
  assign _T_281 = NBufCtr_io_output_count == 3'h1;
  assign _T_287 = io_w_0_en & _T_281;
  assign _T_295 = statesInR_1_io_output_count == 3'h2;
  assign _T_322 = _T_295 ? _T_159 : 7'h0;
  assign _T_331 = _T_330[0];
  assign _T_332 = _T_330[6:1];
  assign _T_358 = _T_295 ? _T_195 : 7'h0;
  assign _T_367 = _T_366[0];
  assign _T_368 = _T_366[6:1];
  assign _T_394 = _T_295 ? _T_231 : 7'h0;
  assign _T_403 = _T_402[0];
  assign _T_404 = _T_402[6:1];
  assign _T_430 = _T_295 ? _T_267 : 7'h0;
  assign _T_440 = _T_438[6:1];
  assign _T_442 = NBufCtr_io_output_count == 3'h2;
  assign _T_448 = io_w_0_en & _T_442;
  assign _T_456 = statesInR_2_io_output_count == 3'h2;
  assign _T_483 = _T_456 ? _T_159 : 7'h0;
  assign _T_492 = _T_491[0];
  assign _T_493 = _T_491[6:1];
  assign _T_519 = _T_456 ? _T_195 : 7'h0;
  assign _T_528 = _T_527[0];
  assign _T_529 = _T_527[6:1];
  assign _T_555 = _T_456 ? _T_231 : 7'h0;
  assign _T_564 = _T_563[0];
  assign _T_565 = _T_563[6:1];
  assign _T_591 = _T_456 ? _T_267 : 7'h0;
  assign _T_601 = _T_599[6:1];
  assign _T_709 = statesOut_2_io_output_count == 3'h0;
  assign _T_712 = statesOut_2_io_output_count == 3'h1;
  assign _T_715 = statesOut_2_io_output_count == 3'h2;
  assign _T_719 = _T_709 ? srams_0_io_output_data_0 : 32'h0;
  assign _T_721 = _T_712 ? srams_1_io_output_data_0 : 32'h0;
  assign _T_723 = _T_715 ? srams_2_io_output_data_0 : 32'h0;
  assign _T_724 = _T_719 | _T_721;
  assign _T_725 = _T_724 | _T_723;
  assign _T_730 = _T_709 ? srams_0_io_output_data_1 : 32'h0;
  assign _T_732 = _T_712 ? srams_1_io_output_data_1 : 32'h0;
  assign _T_734 = _T_715 ? srams_2_io_output_data_1 : 32'h0;
  assign _T_735 = _T_730 | _T_732;
  assign _T_736 = _T_735 | _T_734;
  assign _T_741 = _T_709 ? srams_0_io_output_data_2 : 32'h0;
  assign _T_743 = _T_712 ? srams_1_io_output_data_2 : 32'h0;
  assign _T_745 = _T_715 ? srams_2_io_output_data_2 : 32'h0;
  assign _T_746 = _T_741 | _T_743;
  assign _T_747 = _T_746 | _T_745;
  assign _T_752 = _T_709 ? srams_0_io_output_data_3 : 32'h0;
  assign _T_754 = _T_712 ? srams_1_io_output_data_3 : 32'h0;
  assign _T_756 = _T_715 ? srams_2_io_output_data_3 : 32'h0;
  assign _T_757 = _T_752 | _T_754;
  assign _T_758 = _T_757 | _T_756;
  assign io_output_data_8 = _T_727;
  assign io_output_data_9 = _T_738;
  assign io_output_data_10 = _T_749;
  assign io_output_data_11 = _T_760;
  assign srams_0_io_w_0_addr_0 = _T_124_addr_0;
  assign srams_0_io_w_0_data = _T_124_data;
  assign srams_0_io_w_0_en = _T_124_en;
  assign srams_0_io_r_0_addr_0 = _T_166_addr_0;
  assign srams_0_io_r_0_en = _T_166_en;
  assign srams_0_io_r_1_addr_0 = _T_202_addr_0;
  assign srams_0_io_r_1_en = _T_202_en;
  assign srams_0_io_r_2_addr_0 = _T_238_addr_0;
  assign srams_0_io_r_2_en = _T_238_en;
  assign srams_0_io_r_3_addr_0 = _T_274_addr_0;
  assign srams_0_clock = clock;
  assign srams_1_io_w_0_addr_0 = _T_285_addr_0;
  assign srams_1_io_w_0_data = _T_285_data;
  assign srams_1_io_w_0_en = _T_285_en;
  assign srams_1_io_r_0_addr_0 = _T_327_addr_0;
  assign srams_1_io_r_0_en = _T_327_en;
  assign srams_1_io_r_1_addr_0 = _T_363_addr_0;
  assign srams_1_io_r_1_en = _T_363_en;
  assign srams_1_io_r_2_addr_0 = _T_399_addr_0;
  assign srams_1_io_r_2_en = _T_399_en;
  assign srams_1_io_r_3_addr_0 = _T_435_addr_0;
  assign srams_1_clock = clock;
  assign srams_2_io_w_0_addr_0 = _T_446_addr_0;
  assign srams_2_io_w_0_data = _T_446_data;
  assign srams_2_io_w_0_en = _T_446_en;
  assign srams_2_io_r_0_addr_0 = _T_488_addr_0;
  assign srams_2_io_r_0_en = _T_488_en;
  assign srams_2_io_r_1_addr_0 = _T_524_addr_0;
  assign srams_2_io_r_1_en = _T_524_en;
  assign srams_2_io_r_2_addr_0 = _T_560_addr_0;
  assign srams_2_io_r_2_en = _T_560_en;
  assign srams_2_io_r_3_addr_0 = _T_596_addr_0;
  assign srams_2_clock = clock;
  assign sEn_latch_0_io_input_set = _T_39;
  assign sEn_latch_0_io_input_reset = _T_43;
  assign sEn_latch_0_io_input_asyn_reset = _T_47;
  assign sEn_latch_0_clock = clock;
  assign sEn_latch_0_reset = reset;
  assign sEn_latch_1_io_input_set = _T_57;
  assign sEn_latch_1_io_input_reset = _T_61;
  assign sEn_latch_1_io_input_asyn_reset = _T_65;
  assign sEn_latch_1_clock = clock;
  assign sEn_latch_1_reset = reset;
  assign sEn_latch_2_io_input_set = _T_75;
  assign sEn_latch_2_io_input_reset = _T_79;
  assign sEn_latch_2_io_input_asyn_reset = _T_83;
  assign sEn_latch_2_clock = clock;
  assign sEn_latch_2_reset = reset;
  assign sDone_latch_0_io_input_set = io_sDone_0;
  assign sDone_latch_0_io_input_reset = _T_51;
  assign sDone_latch_0_io_input_asyn_reset = _T_55;
  assign sDone_latch_0_clock = clock;
  assign sDone_latch_0_reset = reset;
  assign sDone_latch_1_io_input_set = io_sDone_1;
  assign sDone_latch_1_io_input_reset = _T_69;
  assign sDone_latch_1_io_input_asyn_reset = _T_73;
  assign sDone_latch_1_clock = clock;
  assign sDone_latch_1_reset = reset;
  assign sDone_latch_2_io_input_set = io_sDone_2;
  assign sDone_latch_2_io_input_reset = _T_87;
  assign sDone_latch_2_io_input_asyn_reset = _T_91;
  assign sDone_latch_2_clock = clock;
  assign sDone_latch_2_reset = reset;
  assign swap = _T_111;
  assign RetimeWrapper_io_flow = 1'h1;
  assign RetimeWrapper_io_in = swap;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_43 = RetimeWrapper_io_out;
  assign RetimeWrapper_1_io_flow = 1'h1;
  assign RetimeWrapper_1_io_in = reset;
  assign RetimeWrapper_1_clock = clock;
  assign RetimeWrapper_1_reset = reset;
  assign _T_47 = RetimeWrapper_1_io_out;
  assign RetimeWrapper_2_io_flow = 1'h1;
  assign RetimeWrapper_2_io_in = swap;
  assign RetimeWrapper_2_clock = clock;
  assign RetimeWrapper_2_reset = reset;
  assign _T_51 = RetimeWrapper_2_io_out;
  assign RetimeWrapper_3_io_flow = 1'h1;
  assign RetimeWrapper_3_io_in = reset;
  assign RetimeWrapper_3_clock = clock;
  assign RetimeWrapper_3_reset = reset;
  assign _T_55 = RetimeWrapper_3_io_out;
  assign RetimeWrapper_4_io_flow = 1'h1;
  assign RetimeWrapper_4_io_in = swap;
  assign RetimeWrapper_4_clock = clock;
  assign RetimeWrapper_4_reset = reset;
  assign _T_61 = RetimeWrapper_4_io_out;
  assign RetimeWrapper_5_io_flow = 1'h1;
  assign RetimeWrapper_5_io_in = reset;
  assign RetimeWrapper_5_clock = clock;
  assign RetimeWrapper_5_reset = reset;
  assign _T_65 = RetimeWrapper_5_io_out;
  assign RetimeWrapper_6_io_flow = 1'h1;
  assign RetimeWrapper_6_io_in = swap;
  assign RetimeWrapper_6_clock = clock;
  assign RetimeWrapper_6_reset = reset;
  assign _T_69 = RetimeWrapper_6_io_out;
  assign RetimeWrapper_7_io_flow = 1'h1;
  assign RetimeWrapper_7_io_in = reset;
  assign RetimeWrapper_7_clock = clock;
  assign RetimeWrapper_7_reset = reset;
  assign _T_73 = RetimeWrapper_7_io_out;
  assign RetimeWrapper_8_io_flow = 1'h1;
  assign RetimeWrapper_8_io_in = swap;
  assign RetimeWrapper_8_clock = clock;
  assign RetimeWrapper_8_reset = reset;
  assign _T_79 = RetimeWrapper_8_io_out;
  assign RetimeWrapper_9_io_flow = 1'h1;
  assign RetimeWrapper_9_io_in = reset;
  assign RetimeWrapper_9_clock = clock;
  assign RetimeWrapper_9_reset = reset;
  assign _T_83 = RetimeWrapper_9_io_out;
  assign RetimeWrapper_10_io_flow = 1'h1;
  assign RetimeWrapper_10_io_in = swap;
  assign RetimeWrapper_10_clock = clock;
  assign RetimeWrapper_10_reset = reset;
  assign _T_87 = RetimeWrapper_10_io_out;
  assign RetimeWrapper_11_io_flow = 1'h1;
  assign RetimeWrapper_11_io_in = reset;
  assign RetimeWrapper_11_clock = clock;
  assign RetimeWrapper_11_reset = reset;
  assign _T_91 = RetimeWrapper_11_io_out;
  assign NBufCtr_io_input_countUp = 1'h0;
  assign NBufCtr_io_input_enable = swap;
  assign NBufCtr_clock = clock;
  assign NBufCtr_reset = reset;
  assign statesInR_0_io_input_countUp = 1'h1;
  assign statesInR_0_io_input_enable = swap;
  assign statesInR_0_clock = clock;
  assign statesInR_0_reset = reset;
  assign statesInR_1_io_input_countUp = 1'h1;
  assign statesInR_1_io_input_enable = swap;
  assign statesInR_1_clock = clock;
  assign statesInR_1_reset = reset;
  assign statesInR_2_io_input_countUp = 1'h1;
  assign statesInR_2_io_input_enable = swap;
  assign statesInR_2_clock = clock;
  assign statesInR_2_reset = reset;
  assign statesOut_0_io_input_countUp = 1'h0;
  assign statesOut_0_io_input_enable = swap;
  assign statesOut_0_clock = clock;
  assign statesOut_0_reset = reset;
  assign statesOut_1_io_input_countUp = 1'h0;
  assign statesOut_1_io_input_enable = swap;
  assign statesOut_1_clock = clock;
  assign statesOut_1_reset = reset;
  assign statesOut_2_io_input_countUp = 1'h0;
  assign statesOut_2_io_input_enable = swap;
  assign statesOut_2_clock = clock;
  assign statesOut_2_reset = reset;
  assign _T_124_addr_0 = io_w_0_addr_0;
  assign _T_124_data = io_w_0_data;
  assign _T_124_en = _T_126;
  assign _T_166_addr_0 = _T_171;
  assign _T_166_en = _T_170;
  assign _T_169 = _T_161;
  assign _T_202_addr_0 = _T_207;
  assign _T_202_en = _T_206;
  assign _T_205 = _T_197;
  assign _T_238_addr_0 = _T_243;
  assign _T_238_en = _T_242;
  assign _T_241 = _T_233;
  assign _T_274_addr_0 = _T_279;
  assign _T_277 = _T_269;
  assign _T_285_addr_0 = io_w_0_addr_0;
  assign _T_285_data = io_w_0_data;
  assign _T_285_en = _T_287;
  assign _T_327_addr_0 = _T_332;
  assign _T_327_en = _T_331;
  assign _T_330 = _T_322;
  assign _T_363_addr_0 = _T_368;
  assign _T_363_en = _T_367;
  assign _T_366 = _T_358;
  assign _T_399_addr_0 = _T_404;
  assign _T_399_en = _T_403;
  assign _T_402 = _T_394;
  assign _T_435_addr_0 = _T_440;
  assign _T_438 = _T_430;
  assign _T_446_addr_0 = io_w_0_addr_0;
  assign _T_446_data = io_w_0_data;
  assign _T_446_en = _T_448;
  assign _T_488_addr_0 = _T_493;
  assign _T_488_en = _T_492;
  assign _T_491 = _T_483;
  assign _T_524_addr_0 = _T_529;
  assign _T_524_en = _T_528;
  assign _T_527 = _T_519;
  assign _T_560_addr_0 = _T_565;
  assign _T_560_en = _T_564;
  assign _T_563 = _T_555;
  assign _T_596_addr_0 = _T_601;
  assign _T_599 = _T_591;
  assign _T_727 = _T_725;
  assign _T_738 = _T_736;
  assign _T_749 = _T_747;
  assign _T_760 = _T_758;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_105 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_105 <= 1'h0;
    end else begin
      _T_105 <= _T_102;
    end
  end
endmodule
module RetimeWrapper_182(
  input        clock,
  input        reset,
  input  [1:0] io_in,
  output [1:0] io_out
);
  wire [1:0] sr_out;
  wire [1:0] sr_in;
  wire  sr_flow;
  wire  sr_reset;
  wire  sr_clock;
  RetimeShiftRegister #(.WIDTH(2), .STAGES(1)) sr (
    .out(sr_out),
    .in(sr_in),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out;
  assign sr_in = io_in;
  assign sr_flow = 1'h1;
  assign sr_reset = reset;
  assign sr_clock = clock;
endmodule
module NBufCtr_36(
  input        clock,
  input        reset,
  input        io_input_countUp,
  input        io_input_enable,
  output [1:0] io_output_count
);
  wire [1:0] _T_8;
  wire [2:0] _T_10;
  wire [1:0] _T_11;
  wire  _T_13;
  wire [1:0] _T_14;
  wire [2:0] _T_16;
  wire [1:0] _T_17;
  wire [1:0] _T_18;
  wire [1:0] _T_19;
  wire [1:0] _T_23;
  wire  _T_25;
  wire [2:0] _T_28;
  wire [2:0] _T_29;
  wire [1:0] _T_30;
  wire [1:0] _T_31;
  wire [1:0] _T_32;
  wire [2:0] _T_34;
  wire [1:0] _T_35;
  wire  _T_37;
  wire [2:0] _T_41;
  wire [1:0] _T_42;
  wire [1:0] _T_43;
  wire [1:0] _T_44;
  wire [2:0] _T_45;
  wire [1:0] _T_46;
  wire [1:0] _T_50;
  wire [1:0] _T_51;
  wire [1:0] _T_54;
  wire [1:0] _T_55;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire [1:0] RetimeWrapper_io_in;
  wire [1:0] RetimeWrapper_io_out;
  wire [1:0] _T_59;
  RetimeWrapper_182 RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_10 = _T_8 + 2'h0;
  assign _T_11 = _T_10[1:0];
  assign _T_13 = _T_11 >= 2'h2;
  assign _T_14 = $signed(_T_8);
  assign _T_16 = $signed(_T_14) + $signed(-2'sh2);
  assign _T_17 = _T_16[1:0];
  assign _T_18 = $signed(_T_17);
  assign _T_19 = $unsigned(_T_18);
  assign _T_23 = _T_13 ? _T_19 : _T_11;
  assign _T_25 = _T_8 == 2'h0;
  assign _T_28 = _T_8 - 2'h1;
  assign _T_29 = $unsigned(_T_28);
  assign _T_30 = _T_29[1:0];
  assign _T_31 = _T_25 ? 2'h1 : _T_30;
  assign _T_32 = io_input_enable ? _T_31 : _T_8;
  assign _T_34 = _T_8 + 2'h1;
  assign _T_35 = _T_34[1:0];
  assign _T_37 = _T_35 >= 2'h2;
  assign _T_41 = $signed(_T_14) + $signed(-2'sh1);
  assign _T_42 = _T_41[1:0];
  assign _T_43 = $signed(_T_42);
  assign _T_44 = $unsigned(_T_43);
  assign _T_45 = 2'h0 + _T_44;
  assign _T_46 = _T_45[1:0];
  assign _T_50 = _T_37 ? _T_46 : _T_35;
  assign _T_51 = io_input_enable ? _T_50 : _T_8;
  assign _T_54 = io_input_countUp ? _T_51 : _T_32;
  assign _T_55 = reset ? 2'h0 : _T_54;
  assign io_output_count = _T_23;
  assign _T_8 = _T_59;
  assign RetimeWrapper_io_in = _T_55;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_59 = RetimeWrapper_io_out;
endmodule
module NBufCtr_38(
  input        clock,
  input        reset,
  input        io_input_countUp,
  input        io_input_enable,
  output [1:0] io_output_count
);
  wire [1:0] _T_8;
  wire [2:0] _T_10;
  wire [1:0] _T_11;
  wire  _T_13;
  wire [1:0] _T_14;
  wire [2:0] _T_16;
  wire [1:0] _T_17;
  wire [1:0] _T_18;
  wire [1:0] _T_19;
  wire [1:0] _T_23;
  wire  _T_25;
  wire [2:0] _T_28;
  wire [2:0] _T_29;
  wire [1:0] _T_30;
  wire [1:0] _T_31;
  wire [1:0] _T_32;
  wire [2:0] _T_45;
  wire [1:0] _T_46;
  wire [1:0] _T_50;
  wire [1:0] _T_51;
  wire [1:0] _T_54;
  wire [1:0] _T_55;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire [1:0] RetimeWrapper_io_in;
  wire [1:0] RetimeWrapper_io_out;
  wire [1:0] _T_59;
  RetimeWrapper_182 RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_10 = _T_8 + 2'h1;
  assign _T_11 = _T_10[1:0];
  assign _T_13 = _T_11 >= 2'h2;
  assign _T_14 = $signed(_T_8);
  assign _T_16 = $signed(_T_14) + $signed(-2'sh1);
  assign _T_17 = _T_16[1:0];
  assign _T_18 = $signed(_T_17);
  assign _T_19 = $unsigned(_T_18);
  assign _T_23 = _T_13 ? _T_19 : _T_11;
  assign _T_25 = _T_8 == 2'h0;
  assign _T_28 = _T_8 - 2'h1;
  assign _T_29 = $unsigned(_T_28);
  assign _T_30 = _T_29[1:0];
  assign _T_31 = _T_25 ? 2'h1 : _T_30;
  assign _T_32 = io_input_enable ? _T_31 : _T_8;
  assign _T_45 = 2'h0 + _T_19;
  assign _T_46 = _T_45[1:0];
  assign _T_50 = _T_13 ? _T_46 : _T_11;
  assign _T_51 = io_input_enable ? _T_50 : _T_8;
  assign _T_54 = io_input_countUp ? _T_51 : _T_32;
  assign _T_55 = reset ? 2'h0 : _T_54;
  assign io_output_count = _T_23;
  assign _T_8 = _T_59;
  assign RetimeWrapper_io_in = _T_55;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_59 = RetimeWrapper_io_out;
endmodule
module NBufSRAMnoBcast_2(
  input         clock,
  input         reset,
  input         io_sEn_0,
  input         io_sEn_1,
  input         io_sDone_0,
  input         io_sDone_1,
  input  [5:0]  io_w_0_addr_0,
  input  [31:0] io_w_0_data,
  input         io_w_0_en,
  input  [5:0]  io_r_0_addr_0,
  input         io_r_0_en,
  input  [5:0]  io_r_1_addr_0,
  input         io_r_1_en,
  input  [5:0]  io_r_2_addr_0,
  input         io_r_2_en,
  input  [5:0]  io_r_3_addr_0,
  input         io_r_3_en,
  output [31:0] io_output_data_4,
  output [31:0] io_output_data_5,
  output [31:0] io_output_data_6,
  output [31:0] io_output_data_7
);
  wire  srams_0_clock;
  wire [5:0] srams_0_io_w_0_addr_0;
  wire [31:0] srams_0_io_w_0_data;
  wire  srams_0_io_w_0_en;
  wire [5:0] srams_0_io_r_0_addr_0;
  wire  srams_0_io_r_0_en;
  wire [5:0] srams_0_io_r_1_addr_0;
  wire  srams_0_io_r_1_en;
  wire [5:0] srams_0_io_r_2_addr_0;
  wire  srams_0_io_r_2_en;
  wire [5:0] srams_0_io_r_3_addr_0;
  wire [31:0] srams_0_io_output_data_0;
  wire [31:0] srams_0_io_output_data_1;
  wire [31:0] srams_0_io_output_data_2;
  wire [31:0] srams_0_io_output_data_3;
  wire  srams_1_clock;
  wire [5:0] srams_1_io_w_0_addr_0;
  wire [31:0] srams_1_io_w_0_data;
  wire  srams_1_io_w_0_en;
  wire [5:0] srams_1_io_r_0_addr_0;
  wire  srams_1_io_r_0_en;
  wire [5:0] srams_1_io_r_1_addr_0;
  wire  srams_1_io_r_1_en;
  wire [5:0] srams_1_io_r_2_addr_0;
  wire  srams_1_io_r_2_en;
  wire [5:0] srams_1_io_r_3_addr_0;
  wire [31:0] srams_1_io_output_data_0;
  wire [31:0] srams_1_io_output_data_1;
  wire [31:0] srams_1_io_output_data_2;
  wire [31:0] srams_1_io_output_data_3;
  wire  sEn_latch_0_clock;
  wire  sEn_latch_0_reset;
  wire  sEn_latch_0_io_input_set;
  wire  sEn_latch_0_io_input_reset;
  wire  sEn_latch_0_io_input_asyn_reset;
  wire  sEn_latch_0_io_output_data;
  wire  sEn_latch_1_clock;
  wire  sEn_latch_1_reset;
  wire  sEn_latch_1_io_input_set;
  wire  sEn_latch_1_io_input_reset;
  wire  sEn_latch_1_io_input_asyn_reset;
  wire  sEn_latch_1_io_output_data;
  wire  sDone_latch_0_clock;
  wire  sDone_latch_0_reset;
  wire  sDone_latch_0_io_input_set;
  wire  sDone_latch_0_io_input_reset;
  wire  sDone_latch_0_io_input_asyn_reset;
  wire  sDone_latch_0_io_output_data;
  wire  sDone_latch_1_clock;
  wire  sDone_latch_1_reset;
  wire  sDone_latch_1_io_input_set;
  wire  sDone_latch_1_io_input_reset;
  wire  sDone_latch_1_io_input_asyn_reset;
  wire  sDone_latch_1_io_output_data;
  wire  swap;
  wire  _T_38;
  wire  _T_39;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire  RetimeWrapper_io_flow;
  wire  RetimeWrapper_io_in;
  wire  RetimeWrapper_io_out;
  wire  _T_43;
  wire  RetimeWrapper_1_clock;
  wire  RetimeWrapper_1_reset;
  wire  RetimeWrapper_1_io_flow;
  wire  RetimeWrapper_1_io_in;
  wire  RetimeWrapper_1_io_out;
  wire  _T_47;
  wire  RetimeWrapper_2_clock;
  wire  RetimeWrapper_2_reset;
  wire  RetimeWrapper_2_io_flow;
  wire  RetimeWrapper_2_io_in;
  wire  RetimeWrapper_2_io_out;
  wire  _T_51;
  wire  RetimeWrapper_3_clock;
  wire  RetimeWrapper_3_reset;
  wire  RetimeWrapper_3_io_flow;
  wire  RetimeWrapper_3_io_in;
  wire  RetimeWrapper_3_io_out;
  wire  _T_55;
  wire  _T_56;
  wire  _T_57;
  wire  RetimeWrapper_4_clock;
  wire  RetimeWrapper_4_reset;
  wire  RetimeWrapper_4_io_flow;
  wire  RetimeWrapper_4_io_in;
  wire  RetimeWrapper_4_io_out;
  wire  _T_61;
  wire  RetimeWrapper_5_clock;
  wire  RetimeWrapper_5_reset;
  wire  RetimeWrapper_5_io_flow;
  wire  RetimeWrapper_5_io_in;
  wire  RetimeWrapper_5_io_out;
  wire  _T_65;
  wire  RetimeWrapper_6_clock;
  wire  RetimeWrapper_6_reset;
  wire  RetimeWrapper_6_io_flow;
  wire  RetimeWrapper_6_io_in;
  wire  RetimeWrapper_6_io_out;
  wire  _T_69;
  wire  RetimeWrapper_7_clock;
  wire  RetimeWrapper_7_reset;
  wire  RetimeWrapper_7_io_flow;
  wire  RetimeWrapper_7_io_in;
  wire  RetimeWrapper_7_io_out;
  wire  _T_73;
  wire  anyEnabled;
  wire  _T_74;
  wire  _T_75;
  wire  _T_76;
  wire  _T_77;
  wire  _T_78;
  wire  _T_79;
  wire  _T_80;
  reg  _T_83;
  reg [31:0] _RAND_0;
  wire  _T_89;
  wire  NBufCtr_clock;
  wire  NBufCtr_reset;
  wire  NBufCtr_io_input_countUp;
  wire  NBufCtr_io_input_enable;
  wire [1:0] NBufCtr_io_output_count;
  wire  statesInR_0_clock;
  wire  statesInR_0_reset;
  wire  statesInR_0_io_input_countUp;
  wire  statesInR_0_io_input_enable;
  wire [1:0] statesInR_0_io_output_count;
  wire  statesInR_1_clock;
  wire  statesInR_1_reset;
  wire  statesInR_1_io_input_countUp;
  wire  statesInR_1_io_input_enable;
  wire [1:0] statesInR_1_io_output_count;
  wire  statesOut_0_clock;
  wire  statesOut_0_reset;
  wire  statesOut_0_io_input_countUp;
  wire  statesOut_0_io_input_enable;
  wire [1:0] statesOut_0_io_output_count;
  wire  statesOut_1_clock;
  wire  statesOut_1_reset;
  wire  statesOut_1_io_input_countUp;
  wire  statesOut_1_io_input_enable;
  wire [1:0] statesOut_1_io_output_count;
  wire  _T_96;
  wire [5:0] _T_100_addr_0;
  wire [31:0] _T_100_data;
  wire  _T_100_en;
  wire  _T_102;
  wire  _T_107;
  wire [6:0] _T_124;
  wire [6:0] _T_126;
  wire [5:0] _T_130_addr_0;
  wire  _T_130_en;
  wire [6:0] _T_133;
  wire  _T_134;
  wire [5:0] _T_135;
  wire [6:0] _T_151;
  wire [6:0] _T_153;
  wire [5:0] _T_157_addr_0;
  wire  _T_157_en;
  wire [6:0] _T_160;
  wire  _T_161;
  wire [5:0] _T_162;
  wire [6:0] _T_178;
  wire [6:0] _T_180;
  wire [5:0] _T_184_addr_0;
  wire  _T_184_en;
  wire [6:0] _T_187;
  wire  _T_188;
  wire [5:0] _T_189;
  wire [6:0] _T_205;
  wire [6:0] _T_207;
  wire [5:0] _T_211_addr_0;
  wire [6:0] _T_214;
  wire [5:0] _T_216;
  wire  _T_218;
  wire [5:0] _T_222_addr_0;
  wire [31:0] _T_222_data;
  wire  _T_222_en;
  wire  _T_224;
  wire  _T_229;
  wire [6:0] _T_248;
  wire [5:0] _T_252_addr_0;
  wire  _T_252_en;
  wire [6:0] _T_255;
  wire  _T_256;
  wire [5:0] _T_257;
  wire [6:0] _T_275;
  wire [5:0] _T_279_addr_0;
  wire  _T_279_en;
  wire [6:0] _T_282;
  wire  _T_283;
  wire [5:0] _T_284;
  wire [6:0] _T_302;
  wire [5:0] _T_306_addr_0;
  wire  _T_306_en;
  wire [6:0] _T_309;
  wire  _T_310;
  wire [5:0] _T_311;
  wire [6:0] _T_329;
  wire [5:0] _T_333_addr_0;
  wire [6:0] _T_336;
  wire [5:0] _T_338;
  wire  _T_378;
  wire  _T_381;
  wire [31:0] _T_385;
  wire [31:0] _T_387;
  wire [31:0] _T_388;
  wire [31:0] _T_390;
  wire [31:0] _T_393;
  wire [31:0] _T_395;
  wire [31:0] _T_396;
  wire [31:0] _T_398;
  wire [31:0] _T_401;
  wire [31:0] _T_403;
  wire [31:0] _T_404;
  wire [31:0] _T_406;
  wire [31:0] _T_409;
  wire [31:0] _T_411;
  wire [31:0] _T_412;
  wire [31:0] _T_414;
  SRAM srams_0 (
    .clock(srams_0_clock),
    .io_w_0_addr_0(srams_0_io_w_0_addr_0),
    .io_w_0_data(srams_0_io_w_0_data),
    .io_w_0_en(srams_0_io_w_0_en),
    .io_r_0_addr_0(srams_0_io_r_0_addr_0),
    .io_r_0_en(srams_0_io_r_0_en),
    .io_r_1_addr_0(srams_0_io_r_1_addr_0),
    .io_r_1_en(srams_0_io_r_1_en),
    .io_r_2_addr_0(srams_0_io_r_2_addr_0),
    .io_r_2_en(srams_0_io_r_2_en),
    .io_r_3_addr_0(srams_0_io_r_3_addr_0),
    .io_output_data_0(srams_0_io_output_data_0),
    .io_output_data_1(srams_0_io_output_data_1),
    .io_output_data_2(srams_0_io_output_data_2),
    .io_output_data_3(srams_0_io_output_data_3)
  );
  SRAM srams_1 (
    .clock(srams_1_clock),
    .io_w_0_addr_0(srams_1_io_w_0_addr_0),
    .io_w_0_data(srams_1_io_w_0_data),
    .io_w_0_en(srams_1_io_w_0_en),
    .io_r_0_addr_0(srams_1_io_r_0_addr_0),
    .io_r_0_en(srams_1_io_r_0_en),
    .io_r_1_addr_0(srams_1_io_r_1_addr_0),
    .io_r_1_en(srams_1_io_r_1_en),
    .io_r_2_addr_0(srams_1_io_r_2_addr_0),
    .io_r_2_en(srams_1_io_r_2_en),
    .io_r_3_addr_0(srams_1_io_r_3_addr_0),
    .io_output_data_0(srams_1_io_output_data_0),
    .io_output_data_1(srams_1_io_output_data_1),
    .io_output_data_2(srams_1_io_output_data_2),
    .io_output_data_3(srams_1_io_output_data_3)
  );
  SRFF sEn_latch_0 (
    .clock(sEn_latch_0_clock),
    .reset(sEn_latch_0_reset),
    .io_input_set(sEn_latch_0_io_input_set),
    .io_input_reset(sEn_latch_0_io_input_reset),
    .io_input_asyn_reset(sEn_latch_0_io_input_asyn_reset),
    .io_output_data(sEn_latch_0_io_output_data)
  );
  SRFF sEn_latch_1 (
    .clock(sEn_latch_1_clock),
    .reset(sEn_latch_1_reset),
    .io_input_set(sEn_latch_1_io_input_set),
    .io_input_reset(sEn_latch_1_io_input_reset),
    .io_input_asyn_reset(sEn_latch_1_io_input_asyn_reset),
    .io_output_data(sEn_latch_1_io_output_data)
  );
  SRFF sDone_latch_0 (
    .clock(sDone_latch_0_clock),
    .reset(sDone_latch_0_reset),
    .io_input_set(sDone_latch_0_io_input_set),
    .io_input_reset(sDone_latch_0_io_input_reset),
    .io_input_asyn_reset(sDone_latch_0_io_input_asyn_reset),
    .io_output_data(sDone_latch_0_io_output_data)
  );
  SRFF sDone_latch_1 (
    .clock(sDone_latch_1_clock),
    .reset(sDone_latch_1_reset),
    .io_input_set(sDone_latch_1_io_input_set),
    .io_input_reset(sDone_latch_1_io_input_reset),
    .io_input_asyn_reset(sDone_latch_1_io_input_asyn_reset),
    .io_output_data(sDone_latch_1_io_output_data)
  );
  RetimeWrapper RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 (
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 (
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 (
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 (
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 (
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 (
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 (
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  NBufCtr_36 NBufCtr (
    .clock(NBufCtr_clock),
    .reset(NBufCtr_reset),
    .io_input_countUp(NBufCtr_io_input_countUp),
    .io_input_enable(NBufCtr_io_input_enable),
    .io_output_count(NBufCtr_io_output_count)
  );
  NBufCtr_36 statesInR_0 (
    .clock(statesInR_0_clock),
    .reset(statesInR_0_reset),
    .io_input_countUp(statesInR_0_io_input_countUp),
    .io_input_enable(statesInR_0_io_input_enable),
    .io_output_count(statesInR_0_io_output_count)
  );
  NBufCtr_38 statesInR_1 (
    .clock(statesInR_1_clock),
    .reset(statesInR_1_reset),
    .io_input_countUp(statesInR_1_io_input_countUp),
    .io_input_enable(statesInR_1_io_input_enable),
    .io_output_count(statesInR_1_io_output_count)
  );
  NBufCtr_36 statesOut_0 (
    .clock(statesOut_0_clock),
    .reset(statesOut_0_reset),
    .io_input_countUp(statesOut_0_io_input_countUp),
    .io_input_enable(statesOut_0_io_input_enable),
    .io_output_count(statesOut_0_io_output_count)
  );
  NBufCtr_38 statesOut_1 (
    .clock(statesOut_1_clock),
    .reset(statesOut_1_reset),
    .io_input_countUp(statesOut_1_io_input_countUp),
    .io_input_enable(statesOut_1_io_input_enable),
    .io_output_count(statesOut_1_io_output_count)
  );
  assign _T_38 = ~ io_sDone_0;
  assign _T_39 = io_sEn_0 & _T_38;
  assign _T_56 = ~ io_sDone_1;
  assign _T_57 = io_sEn_1 & _T_56;
  assign anyEnabled = sEn_latch_0_io_output_data | sEn_latch_1_io_output_data;
  assign _T_74 = sDone_latch_0_io_output_data | io_sDone_0;
  assign _T_75 = sEn_latch_0_io_output_data == _T_74;
  assign _T_76 = sDone_latch_1_io_output_data | io_sDone_1;
  assign _T_77 = sEn_latch_1_io_output_data == _T_76;
  assign _T_78 = _T_75 & _T_77;
  assign _T_79 = _T_78 & anyEnabled;
  assign _T_80 = ~ _T_79;
  assign _T_89 = _T_79 & _T_83;
  assign _T_96 = NBufCtr_io_output_count == 2'h0;
  assign _T_102 = io_w_0_en & _T_96;
  assign _T_107 = statesInR_0_io_output_count == 2'h1;
  assign _T_124 = {io_r_0_addr_0,io_r_0_en};
  assign _T_126 = _T_107 ? _T_124 : 7'h0;
  assign _T_134 = _T_133[0];
  assign _T_135 = _T_133[6:1];
  assign _T_151 = {io_r_1_addr_0,io_r_1_en};
  assign _T_153 = _T_107 ? _T_151 : 7'h0;
  assign _T_161 = _T_160[0];
  assign _T_162 = _T_160[6:1];
  assign _T_178 = {io_r_2_addr_0,io_r_2_en};
  assign _T_180 = _T_107 ? _T_178 : 7'h0;
  assign _T_188 = _T_187[0];
  assign _T_189 = _T_187[6:1];
  assign _T_205 = {io_r_3_addr_0,io_r_3_en};
  assign _T_207 = _T_107 ? _T_205 : 7'h0;
  assign _T_216 = _T_214[6:1];
  assign _T_218 = NBufCtr_io_output_count == 2'h1;
  assign _T_224 = io_w_0_en & _T_218;
  assign _T_229 = statesInR_1_io_output_count == 2'h1;
  assign _T_248 = _T_229 ? _T_124 : 7'h0;
  assign _T_256 = _T_255[0];
  assign _T_257 = _T_255[6:1];
  assign _T_275 = _T_229 ? _T_151 : 7'h0;
  assign _T_283 = _T_282[0];
  assign _T_284 = _T_282[6:1];
  assign _T_302 = _T_229 ? _T_178 : 7'h0;
  assign _T_310 = _T_309[0];
  assign _T_311 = _T_309[6:1];
  assign _T_329 = _T_229 ? _T_205 : 7'h0;
  assign _T_338 = _T_336[6:1];
  assign _T_378 = statesOut_1_io_output_count == 2'h0;
  assign _T_381 = statesOut_1_io_output_count == 2'h1;
  assign _T_385 = _T_378 ? srams_0_io_output_data_0 : 32'h0;
  assign _T_387 = _T_381 ? srams_1_io_output_data_0 : 32'h0;
  assign _T_388 = _T_385 | _T_387;
  assign _T_393 = _T_378 ? srams_0_io_output_data_1 : 32'h0;
  assign _T_395 = _T_381 ? srams_1_io_output_data_1 : 32'h0;
  assign _T_396 = _T_393 | _T_395;
  assign _T_401 = _T_378 ? srams_0_io_output_data_2 : 32'h0;
  assign _T_403 = _T_381 ? srams_1_io_output_data_2 : 32'h0;
  assign _T_404 = _T_401 | _T_403;
  assign _T_409 = _T_378 ? srams_0_io_output_data_3 : 32'h0;
  assign _T_411 = _T_381 ? srams_1_io_output_data_3 : 32'h0;
  assign _T_412 = _T_409 | _T_411;
  assign io_output_data_4 = _T_390;
  assign io_output_data_5 = _T_398;
  assign io_output_data_6 = _T_406;
  assign io_output_data_7 = _T_414;
  assign srams_0_io_w_0_addr_0 = _T_100_addr_0;
  assign srams_0_io_w_0_data = _T_100_data;
  assign srams_0_io_w_0_en = _T_100_en;
  assign srams_0_io_r_0_addr_0 = _T_130_addr_0;
  assign srams_0_io_r_0_en = _T_130_en;
  assign srams_0_io_r_1_addr_0 = _T_157_addr_0;
  assign srams_0_io_r_1_en = _T_157_en;
  assign srams_0_io_r_2_addr_0 = _T_184_addr_0;
  assign srams_0_io_r_2_en = _T_184_en;
  assign srams_0_io_r_3_addr_0 = _T_211_addr_0;
  assign srams_0_clock = clock;
  assign srams_1_io_w_0_addr_0 = _T_222_addr_0;
  assign srams_1_io_w_0_data = _T_222_data;
  assign srams_1_io_w_0_en = _T_222_en;
  assign srams_1_io_r_0_addr_0 = _T_252_addr_0;
  assign srams_1_io_r_0_en = _T_252_en;
  assign srams_1_io_r_1_addr_0 = _T_279_addr_0;
  assign srams_1_io_r_1_en = _T_279_en;
  assign srams_1_io_r_2_addr_0 = _T_306_addr_0;
  assign srams_1_io_r_2_en = _T_306_en;
  assign srams_1_io_r_3_addr_0 = _T_333_addr_0;
  assign srams_1_clock = clock;
  assign sEn_latch_0_io_input_set = _T_39;
  assign sEn_latch_0_io_input_reset = _T_43;
  assign sEn_latch_0_io_input_asyn_reset = _T_47;
  assign sEn_latch_0_clock = clock;
  assign sEn_latch_0_reset = reset;
  assign sEn_latch_1_io_input_set = _T_57;
  assign sEn_latch_1_io_input_reset = _T_61;
  assign sEn_latch_1_io_input_asyn_reset = _T_65;
  assign sEn_latch_1_clock = clock;
  assign sEn_latch_1_reset = reset;
  assign sDone_latch_0_io_input_set = io_sDone_0;
  assign sDone_latch_0_io_input_reset = _T_51;
  assign sDone_latch_0_io_input_asyn_reset = _T_55;
  assign sDone_latch_0_clock = clock;
  assign sDone_latch_0_reset = reset;
  assign sDone_latch_1_io_input_set = io_sDone_1;
  assign sDone_latch_1_io_input_reset = _T_69;
  assign sDone_latch_1_io_input_asyn_reset = _T_73;
  assign sDone_latch_1_clock = clock;
  assign sDone_latch_1_reset = reset;
  assign swap = _T_89;
  assign RetimeWrapper_io_flow = 1'h1;
  assign RetimeWrapper_io_in = swap;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_43 = RetimeWrapper_io_out;
  assign RetimeWrapper_1_io_flow = 1'h1;
  assign RetimeWrapper_1_io_in = reset;
  assign RetimeWrapper_1_clock = clock;
  assign RetimeWrapper_1_reset = reset;
  assign _T_47 = RetimeWrapper_1_io_out;
  assign RetimeWrapper_2_io_flow = 1'h1;
  assign RetimeWrapper_2_io_in = swap;
  assign RetimeWrapper_2_clock = clock;
  assign RetimeWrapper_2_reset = reset;
  assign _T_51 = RetimeWrapper_2_io_out;
  assign RetimeWrapper_3_io_flow = 1'h1;
  assign RetimeWrapper_3_io_in = reset;
  assign RetimeWrapper_3_clock = clock;
  assign RetimeWrapper_3_reset = reset;
  assign _T_55 = RetimeWrapper_3_io_out;
  assign RetimeWrapper_4_io_flow = 1'h1;
  assign RetimeWrapper_4_io_in = swap;
  assign RetimeWrapper_4_clock = clock;
  assign RetimeWrapper_4_reset = reset;
  assign _T_61 = RetimeWrapper_4_io_out;
  assign RetimeWrapper_5_io_flow = 1'h1;
  assign RetimeWrapper_5_io_in = reset;
  assign RetimeWrapper_5_clock = clock;
  assign RetimeWrapper_5_reset = reset;
  assign _T_65 = RetimeWrapper_5_io_out;
  assign RetimeWrapper_6_io_flow = 1'h1;
  assign RetimeWrapper_6_io_in = swap;
  assign RetimeWrapper_6_clock = clock;
  assign RetimeWrapper_6_reset = reset;
  assign _T_69 = RetimeWrapper_6_io_out;
  assign RetimeWrapper_7_io_flow = 1'h1;
  assign RetimeWrapper_7_io_in = reset;
  assign RetimeWrapper_7_clock = clock;
  assign RetimeWrapper_7_reset = reset;
  assign _T_73 = RetimeWrapper_7_io_out;
  assign NBufCtr_io_input_countUp = 1'h0;
  assign NBufCtr_io_input_enable = swap;
  assign NBufCtr_clock = clock;
  assign NBufCtr_reset = reset;
  assign statesInR_0_io_input_countUp = 1'h1;
  assign statesInR_0_io_input_enable = swap;
  assign statesInR_0_clock = clock;
  assign statesInR_0_reset = reset;
  assign statesInR_1_io_input_countUp = 1'h1;
  assign statesInR_1_io_input_enable = swap;
  assign statesInR_1_clock = clock;
  assign statesInR_1_reset = reset;
  assign statesOut_0_io_input_countUp = 1'h0;
  assign statesOut_0_io_input_enable = swap;
  assign statesOut_0_clock = clock;
  assign statesOut_0_reset = reset;
  assign statesOut_1_io_input_countUp = 1'h0;
  assign statesOut_1_io_input_enable = swap;
  assign statesOut_1_clock = clock;
  assign statesOut_1_reset = reset;
  assign _T_100_addr_0 = io_w_0_addr_0;
  assign _T_100_data = io_w_0_data;
  assign _T_100_en = _T_102;
  assign _T_130_addr_0 = _T_135;
  assign _T_130_en = _T_134;
  assign _T_133 = _T_126;
  assign _T_157_addr_0 = _T_162;
  assign _T_157_en = _T_161;
  assign _T_160 = _T_153;
  assign _T_184_addr_0 = _T_189;
  assign _T_184_en = _T_188;
  assign _T_187 = _T_180;
  assign _T_211_addr_0 = _T_216;
  assign _T_214 = _T_207;
  assign _T_222_addr_0 = io_w_0_addr_0;
  assign _T_222_data = io_w_0_data;
  assign _T_222_en = _T_224;
  assign _T_252_addr_0 = _T_257;
  assign _T_252_en = _T_256;
  assign _T_255 = _T_248;
  assign _T_279_addr_0 = _T_284;
  assign _T_279_en = _T_283;
  assign _T_282 = _T_275;
  assign _T_306_addr_0 = _T_311;
  assign _T_306_en = _T_310;
  assign _T_309 = _T_302;
  assign _T_333_addr_0 = _T_338;
  assign _T_336 = _T_329;
  assign _T_390 = _T_388;
  assign _T_398 = _T_396;
  assign _T_406 = _T_404;
  assign _T_414 = _T_412;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_83 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_83 <= 1'h0;
    end else begin
      _T_83 <= _T_80;
    end
  end
endmodule
module FF_30(
  input        clock,
  input        reset,
  input  [1:0] io_input_0_data,
  input        io_input_0_reset,
  output [1:0] io_output_data
);
  reg [1:0] ff;
  reg [31:0] _RAND_0;
  wire [1:0] _T_8;
  wire [1:0] _T_9;
  assign _T_8 = io_input_0_reset ? 2'h1 : io_input_0_data;
  assign _T_9 = io_input_0_reset ? 2'h1 : ff;
  assign io_output_data = _T_9;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  ff = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 2'h1;
    end else begin
      if (io_input_0_reset) begin
        ff <= 2'h1;
      end else begin
        ff <= io_input_0_data;
      end
    end
  end
endmodule
module Parallel(
  input   clock,
  input   reset,
  input   io_input_enable,
  input   io_input_stageDone_0,
  input   io_input_stageDone_1,
  input   io_input_stageMask_0,
  input   io_input_stageMask_1,
  input   io_input_rst,
  output  io_output_done,
  output  io_output_stageEnable_0,
  output  io_output_stageEnable_1,
  output  io_output_rst_en
);
  wire  stateFF_clock;
  wire  stateFF_reset;
  wire [1:0] stateFF_io_input_0_data;
  wire  stateFF_io_input_0_reset;
  wire [1:0] stateFF_io_output_data;
  wire  doneFF_0_clock;
  wire  doneFF_0_reset;
  wire  doneFF_0_io_input_set;
  wire  doneFF_0_io_input_reset;
  wire  doneFF_0_io_input_asyn_reset;
  wire  doneFF_0_io_output_data;
  wire  _T_23;
  wire  _T_24;
  wire  _T_25;
  wire  _T_27;
  wire  _T_29;
  wire  _T_30;
  wire  _T_34;
  wire  _T_40;
  wire  _T_44;
  wire  doneFF_1_clock;
  wire  doneFF_1_reset;
  wire  doneFF_1_io_input_set;
  wire  doneFF_1_io_input_reset;
  wire  doneFF_1_io_input_asyn_reset;
  wire  doneFF_1_io_output_data;
  wire  _T_45;
  wire  _T_46;
  wire  _T_47;
  wire  _T_75;
  wire  _T_77;
  wire  _T_79;
  wire  _T_82;
  wire  _T_84;
  wire  _T_86;
  wire [1:0] _GEN_0;
  wire [1:0] _GEN_1;
  wire  _GEN_2;
  wire  _GEN_3;
  wire [1:0] _GEN_4;
  wire [1:0] _GEN_6;
  wire  _GEN_7;
  wire  _GEN_8;
  wire  _GEN_9;
  wire [1:0] _GEN_10;
  wire  _GEN_11;
  wire  _GEN_12;
  wire  _T_102;
  FF_30 stateFF (
    .clock(stateFF_clock),
    .reset(stateFF_reset),
    .io_input_0_data(stateFF_io_input_0_data),
    .io_input_0_reset(stateFF_io_input_0_reset),
    .io_output_data(stateFF_io_output_data)
  );
  SRFF doneFF_0 (
    .clock(doneFF_0_clock),
    .reset(doneFF_0_reset),
    .io_input_set(doneFF_0_io_input_set),
    .io_input_reset(doneFF_0_io_input_reset),
    .io_input_asyn_reset(doneFF_0_io_input_asyn_reset),
    .io_output_data(doneFF_0_io_output_data)
  );
  SRFF doneFF_1 (
    .clock(doneFF_1_clock),
    .reset(doneFF_1_reset),
    .io_input_set(doneFF_1_io_input_set),
    .io_input_reset(doneFF_1_io_input_reset),
    .io_input_asyn_reset(doneFF_1_io_input_asyn_reset),
    .io_output_data(doneFF_1_io_output_data)
  );
  assign _T_23 = ~ io_input_stageMask_0;
  assign _T_24 = io_input_stageDone_0 | _T_23;
  assign _T_25 = _T_24 & io_input_enable;
  assign _T_27 = stateFF_io_output_data == 2'h3;
  assign _T_29 = stateFF_io_output_data == 2'h1;
  assign _T_30 = _T_27 | _T_29;
  assign _T_34 = _T_30 | _T_27;
  assign _T_40 = _T_30 | io_input_rst;
  assign _T_44 = _T_40 | _T_27;
  assign _T_45 = ~ io_input_stageMask_1;
  assign _T_46 = io_input_stageDone_1 | _T_45;
  assign _T_47 = _T_46 & io_input_enable;
  assign _T_75 = stateFF_io_output_data == 2'h2;
  assign _T_77 = ~ doneFF_0_io_output_data;
  assign _T_79 = io_input_stageMask_0 ? _T_77 : 1'h0;
  assign _T_82 = ~ doneFF_1_io_output_data;
  assign _T_84 = io_input_stageMask_1 ? _T_82 : 1'h0;
  assign _T_86 = doneFF_0_io_output_data & doneFF_1_io_output_data;
  assign _GEN_0 = _T_86 ? 2'h3 : stateFF_io_output_data;
  assign _GEN_1 = _T_27 ? 2'h1 : stateFF_io_output_data;
  assign _GEN_2 = _T_75 ? _T_79 : 1'h0;
  assign _GEN_3 = _T_75 ? _T_84 : 1'h0;
  assign _GEN_4 = _T_75 ? _GEN_0 : _GEN_1;
  assign _GEN_6 = _T_29 ? 2'h2 : _GEN_4;
  assign _GEN_7 = _T_29 ? 1'h0 : _GEN_2;
  assign _GEN_8 = _T_29 ? 1'h0 : _GEN_3;
  assign _GEN_9 = io_input_enable ? _T_29 : 1'h0;
  assign _GEN_10 = io_input_enable ? _GEN_6 : 2'h1;
  assign _GEN_11 = io_input_enable ? _GEN_7 : 1'h0;
  assign _GEN_12 = io_input_enable ? _GEN_8 : 1'h0;
  assign _T_102 = _T_75 & _T_86;
  assign io_output_done = _T_102;
  assign io_output_stageEnable_0 = _GEN_11;
  assign io_output_stageEnable_1 = _GEN_12;
  assign io_output_rst_en = _GEN_9;
  assign stateFF_io_input_0_data = _GEN_10;
  assign stateFF_io_input_0_reset = io_input_rst;
  assign stateFF_clock = clock;
  assign stateFF_reset = reset;
  assign doneFF_0_io_input_set = _T_25;
  assign doneFF_0_io_input_reset = _T_44;
  assign doneFF_0_io_input_asyn_reset = _T_34;
  assign doneFF_0_clock = clock;
  assign doneFF_0_reset = reset;
  assign doneFF_1_io_input_set = _T_47;
  assign doneFF_1_io_input_reset = _T_44;
  assign doneFF_1_io_input_asyn_reset = _T_34;
  assign doneFF_1_clock = clock;
  assign doneFF_1_reset = reset;
endmodule
module Innerpipe(
  input   clock,
  input   reset,
  input   io_input_enable,
  input   io_input_ctr_done,
  input   io_input_rst,
  output  io_output_done,
  output  io_output_ctr_inc
);
  wire  SRFF_clock;
  wire  SRFF_reset;
  wire  SRFF_io_input_set;
  wire  SRFF_io_input_reset;
  wire  SRFF_io_input_asyn_reset;
  wire  SRFF_io_output_data;
  wire  FF_clock;
  wire  FF_reset;
  wire [31:0] FF_io_input_0_data;
  wire [31:0] FF_io_input_0_init;
  wire  FF_io_input_0_enable;
  wire  FF_io_input_0_reset;
  wire [31:0] FF_io_output_data;
  wire  _T_19;
  wire  _T_20;
  wire  _T_22;
  wire  _T_24;
  wire  _T_25;
  wire  _T_26;
  wire  _T_28;
  wire  _T_31;
  wire  _T_32;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire  RetimeWrapper_io_flow;
  wire  RetimeWrapper_io_in;
  wire  RetimeWrapper_io_out;
  wire  _T_39;
  wire [1:0] _T_45;
  wire [1:0] _T_48;
  wire [1:0] _GEN_0;
  wire  _T_50;
  wire  _T_53;
  wire  RetimeWrapper_1_clock;
  wire  RetimeWrapper_1_reset;
  wire  RetimeWrapper_1_io_flow;
  wire  RetimeWrapper_1_io_in;
  wire  RetimeWrapper_1_io_out;
  wire  _T_57;
  wire  _T_58;
  wire  _T_59;
  wire  _T_60;
  wire  _GEN_3;
  wire  _T_76;
  wire  _T_84;
  wire [32:0] _T_92;
  wire [31:0] _T_93;
  wire [31:0] _T_94;
  wire [31:0] _GEN_9;
  wire  _GEN_10;
  wire  _GEN_11;
  wire [31:0] _GEN_13;
  wire  _GEN_14;
  wire  _GEN_16;
  wire [31:0] _GEN_17;
  wire  _T_97;
  wire  _T_98;
  wire  _GEN_18;
  wire  _GEN_20;
  wire [31:0] _GEN_21;
  SRFF SRFF (
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output_data(SRFF_io_output_data)
  );
  FF_1 FF (
    .clock(FF_clock),
    .reset(FF_reset),
    .io_input_0_data(FF_io_input_0_data),
    .io_input_0_init(FF_io_input_0_init),
    .io_input_0_enable(FF_io_input_0_enable),
    .io_input_0_reset(FF_io_input_0_reset),
    .io_output_data(FF_io_output_data)
  );
  RetimeWrapper RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 (
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign _T_19 = ~ io_input_enable;
  assign _T_20 = _T_19 | io_input_rst;
  assign _T_22 = FF_io_output_data != 32'h3;
  assign _T_24 = FF_io_output_data != 32'h1;
  assign _T_25 = _T_22 & _T_24;
  assign _T_26 = _T_20 | _T_25;
  assign _T_28 = FF_io_output_data != 32'h2;
  assign _T_31 = _T_28 & _T_24;
  assign _T_32 = _T_31 | SRFF_io_output_data;
  assign _T_39 = FF_io_output_data == 32'h1;
  assign _T_45 = io_input_ctr_done ? 2'h3 : 2'h2;
  assign _T_48 = io_input_ctr_done ? 2'h3 : 2'h1;
  assign _GEN_0 = _T_26 ? _T_48 : _T_45;
  assign _T_50 = FF_io_output_data == 32'h2;
  assign _T_53 = _T_28 | SRFF_io_output_data;
  assign _T_58 = _T_57 | io_input_rst;
  assign _T_59 = ~ _T_58;
  assign _T_60 = io_input_enable & _T_59;
  assign _GEN_3 = io_input_ctr_done ? 1'h0 : _T_60;
  assign _T_76 = FF_io_output_data == 32'h3;
  assign _T_84 = FF_io_output_data >= 32'h4;
  assign _T_92 = FF_io_output_data + 32'h1;
  assign _T_93 = _T_92[31:0];
  assign _T_94 = _T_84 ? 32'h2 : _T_93;
  assign _GEN_9 = _T_76 ? 32'h2 : _T_94;
  assign _GEN_10 = _T_50 ? _GEN_3 : 1'h0;
  assign _GEN_11 = _T_50 ? io_input_ctr_done : 1'h0;
  assign _GEN_13 = _T_50 ? {{30'd0}, _T_45} : _GEN_9;
  assign _GEN_14 = _T_39 ? 1'h0 : _GEN_11;
  assign _GEN_16 = _T_39 ? 1'h0 : _GEN_10;
  assign _GEN_17 = _T_39 ? {{30'd0}, _GEN_0} : _GEN_13;
  assign _T_97 = _T_50 & io_input_ctr_done;
  assign _T_98 = io_input_ctr_done | _T_97;
  assign _GEN_18 = io_input_enable ? _GEN_14 : _T_98;
  assign _GEN_20 = io_input_enable ? _GEN_16 : 1'h0;
  assign _GEN_21 = io_input_enable ? _GEN_17 : 32'h2;
  assign io_output_done = _GEN_18;
  assign io_output_ctr_inc = _GEN_20;
  assign SRFF_io_input_set = io_input_rst;
  assign SRFF_io_input_reset = io_input_enable;
  assign SRFF_io_input_asyn_reset = io_input_enable;
  assign SRFF_clock = clock;
  assign SRFF_reset = reset;
  assign FF_io_input_0_data = _GEN_21;
  assign FF_io_input_0_init = 32'h2;
  assign FF_io_input_0_enable = 1'h1;
  assign FF_io_input_0_reset = 1'h0;
  assign FF_clock = clock;
  assign FF_reset = reset;
  assign RetimeWrapper_io_flow = 1'h1;
  assign RetimeWrapper_io_in = _T_32;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign RetimeWrapper_1_io_flow = 1'h1;
  assign RetimeWrapper_1_io_in = _T_53;
  assign RetimeWrapper_1_clock = clock;
  assign RetimeWrapper_1_reset = reset;
  assign _T_57 = RetimeWrapper_1_io_out;
endmodule
module FF_35(
  input        clock,
  input        reset,
  input  [5:0] io_input_0_data,
  input        io_input_0_enable,
  input        io_input_0_reset,
  output [5:0] io_output_data
);
  reg [5:0] ff;
  reg [31:0] _RAND_0;
  wire [5:0] _T_7;
  wire [5:0] _T_8;
  wire [5:0] _T_9;
  assign _T_7 = io_input_0_enable ? io_input_0_data : ff;
  assign _T_8 = io_input_0_reset ? 6'h0 : _T_7;
  assign _T_9 = io_input_0_reset ? 6'h0 : ff;
  assign io_output_data = _T_9;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  ff = _RAND_0[5:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 6'h0;
    end else begin
      if (io_input_0_reset) begin
        ff <= 6'h0;
      end else begin
        if (io_input_0_enable) begin
          ff <= io_input_0_data;
        end
      end
    end
  end
endmodule
module CompactingCounter(
  input        clock,
  input        reset,
  input        io_input_reset,
  input        io_input_enables_0,
  output [5:0] io_output_count
);
  wire  base_clock;
  wire  base_reset;
  wire [5:0] base_io_input_0_data;
  wire  base_io_input_0_enable;
  wire  base_io_input_0_reset;
  wire [5:0] base_io_output_data;
  wire [5:0] count;
  wire [5:0] num_enabled;
  wire [6:0] _T_17;
  wire [5:0] _T_18;
  wire [5:0] newval;
  wire  isMax;
  wire [6:0] _T_24;
  wire [5:0] _T_25;
  wire [5:0] _T_26;
  wire [5:0] next;
  wire [5:0] _T_28;
  wire [5:0] _T_29;
  FF_35 base (
    .clock(base_clock),
    .reset(base_reset),
    .io_input_0_data(base_io_input_0_data),
    .io_input_0_enable(base_io_input_0_enable),
    .io_input_0_reset(base_io_input_0_reset),
    .io_output_data(base_io_output_data)
  );
  assign count = $signed(base_io_output_data);
  assign num_enabled = io_input_enables_0 ? $signed(6'sh1) : $signed(6'sh0);
  assign _T_17 = $signed(count) + $signed(num_enabled);
  assign _T_18 = _T_17[5:0];
  assign newval = $signed(_T_18);
  assign isMax = $signed(newval) >= $signed(6'sh10);
  assign _T_24 = $signed(newval) - $signed(6'sh10);
  assign _T_25 = _T_24[5:0];
  assign _T_26 = $signed(_T_25);
  assign next = isMax ? $signed(_T_26) : $signed(newval);
  assign _T_28 = $unsigned(next);
  assign _T_29 = io_input_reset ? 6'h0 : _T_28;
  assign io_output_count = count;
  assign base_io_input_0_data = _T_29;
  assign base_io_input_0_enable = io_input_enables_0;
  assign base_io_input_0_reset = io_input_reset;
  assign base_clock = clock;
  assign base_reset = reset;
endmodule
module CompactingIncDincCtr(
  input   clock,
  input   reset,
  input   io_input_inc_en_0,
  input   io_input_dinc_en_0,
  output  io_output_empty,
  output  io_output_full
);
  reg [31:0] cnt;
  reg [31:0] _RAND_0;
  wire [5:0] numPushed;
  wire [5:0] numPopped;
  wire [31:0] _GEN_0;
  wire [32:0] _T_21;
  wire [31:0] _T_22;
  wire [31:0] _T_23;
  wire [31:0] _GEN_1;
  wire [32:0] _T_24;
  wire [31:0] _T_25;
  wire [31:0] _T_26;
  wire  _T_32;
  wire  _T_40;
  assign numPushed = io_input_inc_en_0 ? $signed(6'sh1) : $signed(6'sh0);
  assign numPopped = io_input_dinc_en_0 ? $signed(6'sh1) : $signed(6'sh0);
  assign _GEN_0 = {{26{numPushed[5]}},numPushed};
  assign _T_21 = $signed(cnt) + $signed(_GEN_0);
  assign _T_22 = _T_21[31:0];
  assign _T_23 = $signed(_T_22);
  assign _GEN_1 = {{26{numPopped[5]}},numPopped};
  assign _T_24 = $signed(_T_23) - $signed(_GEN_1);
  assign _T_25 = _T_24[31:0];
  assign _T_26 = $signed(_T_25);
  assign _T_32 = $signed(cnt) == $signed(32'sh0);
  assign _T_40 = $signed(cnt) == $signed(32'sh10);
  assign io_output_empty = _T_32;
  assign io_output_full = _T_40;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  cnt = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      cnt <= 32'sh0;
    end else begin
      cnt <= _T_26;
    end
  end
endmodule
module Mem1D_40(
  input         clock,
  input  [3:0]  io_w_addr,
  input  [95:0] io_w_data,
  input         io_w_en,
  input  [3:0]  io_r_addr,
  output [95:0] io_output_data
);
  reg [95:0] _T_14 [0:15];
  reg [95:0] _RAND_0;
  wire [95:0] _T_14__T_17_data;
  wire [3:0] _T_14__T_17_addr;
  wire [95:0] _T_14__T_16_data;
  wire [3:0] _T_14__T_16_addr;
  wire  _T_14__T_16_mask;
  wire  _T_14__T_16_en;
  assign _T_14__T_17_addr = io_r_addr;
  assign _T_14__T_17_data = _T_14[_T_14__T_17_addr];
  assign _T_14__T_16_data = io_w_data;
  assign _T_14__T_16_addr = io_w_addr;
  assign _T_14__T_16_mask = io_w_en;
  assign _T_14__T_16_en = io_w_en;
  assign io_output_data = _T_14__T_17_data;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {3{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    _T_14[initvar] = _RAND_0[95:0];
  `endif // RANDOMIZE_MEM_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(_T_14__T_16_en & _T_14__T_16_mask) begin
      _T_14[_T_14__T_16_addr] <= _T_14__T_16_data;
    end
  end
endmodule
module Compactor(
  input  [95:0] io_in_0_data,
  output [95:0] io_out_0_data
);
  assign io_out_0_data = io_in_0_data;
endmodule
module CompactingEnqNetwork(
  input  [5:0]  io_headCnt,
  input  [95:0] io_in_0_data,
  input         io_in_0_en,
  output [95:0] io_out_0_data,
  output        io_out_0_en
);
  wire [5:0] numEnabled;
  wire [95:0] compactor_io_in_0_data;
  wire [95:0] compactor_io_out_0_data;
  wire [5:0] _GEN_0;
  wire [5:0] current_base_bank;
  wire [5:0] _T_14;
  wire [6:0] _T_15;
  wire [5:0] _T_16;
  wire [5:0] _T_17;
  wire [6:0] _T_19;
  wire [5:0] _T_20;
  wire [5:0] upper;
  wire  _T_22;
  wire [5:0] num_straddling;
  wire [6:0] _T_25;
  wire [5:0] _T_26;
  wire [5:0] num_straight;
  wire  _T_28;
  wire  _T_30;
  wire  _T_36;
  wire  _T_37;
  wire  _T_38;
  wire [6:0] _T_45;
  wire [5:0] _T_46;
  wire [5:0] _T_47;
  wire [6:0] _T_49;
  wire [5:0] _T_50;
  wire [5:0] _T_51;
  wire [5:0] _T_52;
  wire [5:0] _T_54;
  wire  _T_56;
  wire [95:0] _T_57;
  Compactor compactor (
    .io_in_0_data(compactor_io_in_0_data),
    .io_out_0_data(compactor_io_out_0_data)
  );
  assign numEnabled = io_in_0_en ? 6'h1 : 6'h0;
  assign _GEN_0 = $signed(io_headCnt) % $signed(6'sh1);
  assign current_base_bank = _GEN_0[5:0];
  assign _T_14 = $signed(numEnabled);
  assign _T_15 = $signed(current_base_bank) + $signed(_T_14);
  assign _T_16 = _T_15[5:0];
  assign _T_17 = $signed(_T_16);
  assign _T_19 = $signed(_T_17) - $signed(6'sh1);
  assign _T_20 = _T_19[5:0];
  assign upper = $signed(_T_20);
  assign _T_22 = $signed(upper) < $signed(6'sh0);
  assign num_straddling = _T_22 ? $signed(6'sh0) : $signed(upper);
  assign _T_25 = $signed(_T_14) - $signed(num_straddling);
  assign _T_26 = _T_25[5:0];
  assign num_straight = $signed(_T_26);
  assign _T_28 = $signed(6'sh0) < $signed(num_straddling);
  assign _T_30 = $signed(6'sh0) >= $signed(current_base_bank);
  assign _T_36 = $signed(6'sh0) < $signed(_T_17);
  assign _T_37 = _T_30 & _T_36;
  assign _T_38 = _T_28 | _T_37;
  assign _T_45 = $signed(6'sh0) + $signed(num_straight);
  assign _T_46 = _T_45[5:0];
  assign _T_47 = $signed(_T_46);
  assign _T_49 = $signed(6'sh0) - $signed(current_base_bank);
  assign _T_50 = _T_49[5:0];
  assign _T_51 = $signed(_T_50);
  assign _T_52 = _T_28 ? $signed(_T_47) : $signed(_T_51);
  assign _T_54 = $unsigned(_T_52);
  assign _T_56 = 6'h0 == _T_54;
  assign _T_57 = _T_56 ? compactor_io_out_0_data : 96'h0;
  assign io_out_0_data = _T_57;
  assign io_out_0_en = _T_38;
  assign compactor_io_in_0_data = io_in_0_data;
endmodule
module CompactingDeqNetwork(
  input  [5:0]  io_tailCnt,
  input  [95:0] io_input_data_0,
  output [95:0] io_output_data_0
);
  wire [5:0] _GEN_0;
  wire [5:0] current_base_bank;
  wire [5:0] _T_42;
  wire [6:0] _T_43;
  wire [5:0] _T_44;
  wire [5:0] _GEN_1;
  wire [5:0] _T_46;
  wire  _T_49;
  wire [95:0] _T_50;
  assign _GEN_0 = $signed(io_tailCnt) % $signed(6'sh1);
  assign current_base_bank = _GEN_0[5:0];
  assign _T_42 = $unsigned(current_base_bank);
  assign _T_43 = _T_42 + 6'h0;
  assign _T_44 = _T_43[5:0];
  assign _GEN_1 = _T_44 % 6'h1;
  assign _T_46 = _GEN_1[5:0];
  assign _T_49 = 6'h0 == _T_46;
  assign _T_50 = _T_49 ? io_input_data_0 : 96'h0;
  assign io_output_data_0 = _T_50;
endmodule
module GeneralFIFO(
  input         clock,
  input         reset,
  input  [95:0] io_in_0_data,
  input         io_in_0_en,
  output [95:0] io_out_0,
  input         io_deq_0,
  output        io_empty,
  output        io_full
);
  wire  headCtr_clock;
  wire  headCtr_reset;
  wire  headCtr_io_input_reset;
  wire  headCtr_io_input_enables_0;
  wire [5:0] headCtr_io_output_count;
  wire  tailCtr_clock;
  wire  tailCtr_reset;
  wire  tailCtr_io_input_reset;
  wire  tailCtr_io_input_enables_0;
  wire [5:0] tailCtr_io_output_count;
  wire  elements_clock;
  wire  elements_reset;
  wire  elements_io_input_inc_en_0;
  wire  elements_io_input_dinc_en_0;
  wire  elements_io_output_empty;
  wire  elements_io_output_full;
  wire  m_0_clock;
  wire [3:0] m_0_io_w_addr;
  wire [95:0] m_0_io_w_data;
  wire  m_0_io_w_en;
  wire [3:0] m_0_io_r_addr;
  wire [95:0] m_0_io_output_data;
  wire [5:0] enqCompactor_io_headCnt;
  wire [95:0] enqCompactor_io_in_0_data;
  wire  enqCompactor_io_in_0_en;
  wire [95:0] enqCompactor_io_out_0_data;
  wire  enqCompactor_io_out_0_en;
  wire [5:0] _GEN_0;
  wire [5:0] active_w_bank;
  wire [6:0] active_w_addr;
  wire  _T_24;
  wire [7:0] _T_26;
  wire [6:0] _T_27;
  wire [6:0] _T_28;
  wire [6:0] _T_29;
  wire [6:0] _T_30;
  wire [5:0] deqCompactor_io_tailCnt;
  wire [95:0] deqCompactor_io_input_data_0;
  wire [95:0] deqCompactor_io_output_data_0;
  wire [5:0] _GEN_1;
  wire [5:0] active_r_bank;
  wire [6:0] active_r_addr;
  wire  _T_34;
  wire [7:0] _T_36;
  wire [6:0] _T_37;
  wire [6:0] _T_38;
  wire [6:0] _T_39;
  wire [6:0] _T_40;
  CompactingCounter headCtr (
    .clock(headCtr_clock),
    .reset(headCtr_reset),
    .io_input_reset(headCtr_io_input_reset),
    .io_input_enables_0(headCtr_io_input_enables_0),
    .io_output_count(headCtr_io_output_count)
  );
  CompactingCounter tailCtr (
    .clock(tailCtr_clock),
    .reset(tailCtr_reset),
    .io_input_reset(tailCtr_io_input_reset),
    .io_input_enables_0(tailCtr_io_input_enables_0),
    .io_output_count(tailCtr_io_output_count)
  );
  CompactingIncDincCtr elements (
    .clock(elements_clock),
    .reset(elements_reset),
    .io_input_inc_en_0(elements_io_input_inc_en_0),
    .io_input_dinc_en_0(elements_io_input_dinc_en_0),
    .io_output_empty(elements_io_output_empty),
    .io_output_full(elements_io_output_full)
  );
  Mem1D_40 m_0 (
    .clock(m_0_clock),
    .io_w_addr(m_0_io_w_addr),
    .io_w_data(m_0_io_w_data),
    .io_w_en(m_0_io_w_en),
    .io_r_addr(m_0_io_r_addr),
    .io_output_data(m_0_io_output_data)
  );
  CompactingEnqNetwork enqCompactor (
    .io_headCnt(enqCompactor_io_headCnt),
    .io_in_0_data(enqCompactor_io_in_0_data),
    .io_in_0_en(enqCompactor_io_in_0_en),
    .io_out_0_data(enqCompactor_io_out_0_data),
    .io_out_0_en(enqCompactor_io_out_0_en)
  );
  CompactingDeqNetwork deqCompactor (
    .io_tailCnt(deqCompactor_io_tailCnt),
    .io_input_data_0(deqCompactor_io_input_data_0),
    .io_output_data_0(deqCompactor_io_output_data_0)
  );
  assign _GEN_0 = $signed(headCtr_io_output_count) % $signed(6'sh1);
  assign active_w_bank = _GEN_0[5:0];
  assign active_w_addr = $signed(headCtr_io_output_count) / $signed(6'sh1);
  assign _T_24 = $signed(6'sh0) < $signed(active_w_bank);
  assign _T_26 = $signed(active_w_addr) + $signed(7'sh1);
  assign _T_27 = _T_26[6:0];
  assign _T_28 = $signed(_T_27);
  assign _T_29 = _T_24 ? $signed(_T_28) : $signed(active_w_addr);
  assign _T_30 = $unsigned(_T_29);
  assign _GEN_1 = $signed(tailCtr_io_output_count) % $signed(6'sh1);
  assign active_r_bank = _GEN_1[5:0];
  assign active_r_addr = $signed(tailCtr_io_output_count) / $signed(6'sh1);
  assign _T_34 = $signed(6'sh0) < $signed(active_r_bank);
  assign _T_36 = $signed(active_r_addr) + $signed(7'sh1);
  assign _T_37 = _T_36[6:0];
  assign _T_38 = $signed(_T_37);
  assign _T_39 = _T_34 ? $signed(_T_38) : $signed(active_r_addr);
  assign _T_40 = $unsigned(_T_39);
  assign io_out_0 = deqCompactor_io_output_data_0;
  assign io_empty = elements_io_output_empty;
  assign io_full = elements_io_output_full;
  assign headCtr_io_input_reset = reset;
  assign headCtr_io_input_enables_0 = io_in_0_en;
  assign headCtr_clock = clock;
  assign headCtr_reset = reset;
  assign tailCtr_io_input_reset = reset;
  assign tailCtr_io_input_enables_0 = io_deq_0;
  assign tailCtr_clock = clock;
  assign tailCtr_reset = reset;
  assign elements_io_input_inc_en_0 = io_in_0_en;
  assign elements_io_input_dinc_en_0 = io_deq_0;
  assign elements_clock = clock;
  assign elements_reset = reset;
  assign m_0_io_w_addr = _T_30[3:0];
  assign m_0_io_w_data = enqCompactor_io_out_0_data;
  assign m_0_io_w_en = enqCompactor_io_out_0_en;
  assign m_0_io_r_addr = _T_40[3:0];
  assign m_0_clock = clock;
  assign enqCompactor_io_headCnt = headCtr_io_output_count;
  assign enqCompactor_io_in_0_data = io_in_0_data;
  assign enqCompactor_io_in_0_en = io_in_0_en;
  assign deqCompactor_io_tailCnt = tailCtr_io_output_count;
  assign deqCompactor_io_input_data_0 = m_0_io_output_data;
endmodule
module Counter_1(
  input         clock,
  input         reset,
  input  [31:0] io_input_stops_0,
  input         io_input_reset,
  input         io_input_enable,
  output [31:0] io_output_counts_0,
  output        io_output_done
);
  wire  ctrs_0_clock;
  wire  ctrs_0_reset;
  wire [31:0] ctrs_0_io_input_stop;
  wire [31:0] ctrs_0_io_input_stride;
  wire  ctrs_0_io_input_reset;
  wire  ctrs_0_io_input_enable;
  wire  ctrs_0_io_input_saturate;
  wire [31:0] ctrs_0_io_output_count_0;
  wire  ctrs_0_io_output_done;
  reg  wasDone;
  reg [31:0] _RAND_0;
  wire  _T_29;
  wire  _T_30;
  wire  _T_31;
  SingleCounter_1 ctrs_0 (
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_input_stop(ctrs_0_io_input_stop),
    .io_input_stride(ctrs_0_io_input_stride),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_input_saturate(ctrs_0_io_input_saturate),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_done(ctrs_0_io_output_done)
  );
  assign _T_29 = io_input_enable & ctrs_0_io_output_done;
  assign _T_30 = ~ wasDone;
  assign _T_31 = _T_29 & _T_30;
  assign io_output_counts_0 = ctrs_0_io_output_count_0;
  assign io_output_done = _T_31;
  assign ctrs_0_io_input_stop = io_input_stops_0;
  assign ctrs_0_io_input_stride = 32'sh1;
  assign ctrs_0_io_input_reset = io_input_reset;
  assign ctrs_0_io_input_enable = io_input_enable;
  assign ctrs_0_io_input_saturate = 1'h0;
  assign ctrs_0_clock = clock;
  assign ctrs_0_reset = reset;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= ctrs_0_io_output_done;
    end
  end
endmodule
module Streaminner(
  input   io_input_ctr_done,
  output  io_output_done
);
  assign io_output_done = io_input_ctr_done;
endmodule
module NBufCtr_46(
  input        clock,
  input        reset,
  input        io_input_enable,
  output [1:0] io_output_count
);
  wire [1:0] _T_8;
  wire [2:0] _T_9;
  wire [1:0] _T_10;
  wire  _T_12;
  wire [2:0] _T_16;
  wire [2:0] _T_17;
  wire [1:0] _T_18;
  wire [1:0] _T_21;
  wire  _T_23;
  wire [2:0] _T_26;
  wire [2:0] _T_27;
  wire [1:0] _T_28;
  wire [1:0] _T_29;
  wire [1:0] _T_30;
  wire [1:0] _T_54;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire [1:0] RetimeWrapper_io_in;
  wire [1:0] RetimeWrapper_io_out;
  wire [1:0] _T_58;
  RetimeWrapper_182 RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_9 = _T_8 + 2'h0;
  assign _T_10 = _T_9[1:0];
  assign _T_12 = _T_10 >= 2'h2;
  assign _T_16 = _T_10 - 2'h2;
  assign _T_17 = $unsigned(_T_16);
  assign _T_18 = _T_17[1:0];
  assign _T_21 = _T_12 ? _T_18 : _T_10;
  assign _T_23 = _T_8 == 2'h0;
  assign _T_26 = _T_8 - 2'h1;
  assign _T_27 = $unsigned(_T_26);
  assign _T_28 = _T_27[1:0];
  assign _T_29 = _T_23 ? 2'h1 : _T_28;
  assign _T_30 = io_input_enable ? _T_29 : _T_8;
  assign _T_54 = reset ? 2'h0 : _T_30;
  assign io_output_count = _T_21;
  assign _T_8 = _T_58;
  assign RetimeWrapper_io_in = _T_54;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_58 = RetimeWrapper_io_out;
endmodule
module NBufFF_4(
  input         clock,
  input         reset,
  input         io_sEn_0,
  input         io_sEn_1,
  input         io_sDone_0,
  input         io_sDone_1,
  input  [31:0] io_input_0_data,
  input         io_input_0_enable,
  input         io_input_0_reset,
  output [31:0] io_output_1_data
);
  wire  ff_0_clock;
  wire  ff_0_reset;
  wire [31:0] ff_0_io_input_0_data;
  wire [31:0] ff_0_io_input_0_init;
  wire  ff_0_io_input_0_enable;
  wire  ff_0_io_input_0_reset;
  wire [31:0] ff_0_io_output_data;
  wire  ff_1_clock;
  wire  ff_1_reset;
  wire [31:0] ff_1_io_input_0_data;
  wire [31:0] ff_1_io_input_0_init;
  wire  ff_1_io_input_0_enable;
  wire  ff_1_io_input_0_reset;
  wire [31:0] ff_1_io_output_data;
  wire  sEn_latch_0_clock;
  wire  sEn_latch_0_reset;
  wire  sEn_latch_0_io_input_set;
  wire  sEn_latch_0_io_input_reset;
  wire  sEn_latch_0_io_input_asyn_reset;
  wire  sEn_latch_0_io_output_data;
  wire  sEn_latch_1_clock;
  wire  sEn_latch_1_reset;
  wire  sEn_latch_1_io_input_set;
  wire  sEn_latch_1_io_input_reset;
  wire  sEn_latch_1_io_input_asyn_reset;
  wire  sEn_latch_1_io_output_data;
  wire  sDone_latch_0_clock;
  wire  sDone_latch_0_reset;
  wire  sDone_latch_0_io_input_set;
  wire  sDone_latch_0_io_input_reset;
  wire  sDone_latch_0_io_input_asyn_reset;
  wire  sDone_latch_0_io_output_data;
  wire  sDone_latch_1_clock;
  wire  sDone_latch_1_reset;
  wire  sDone_latch_1_io_input_set;
  wire  sDone_latch_1_io_input_reset;
  wire  sDone_latch_1_io_input_asyn_reset;
  wire  sDone_latch_1_io_output_data;
  wire  swap;
  wire  _T_20;
  wire  _T_21;
  wire  _T_22;
  wire  _T_23;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire  RetimeWrapper_io_flow;
  wire  RetimeWrapper_io_in;
  wire  RetimeWrapper_io_out;
  wire  _T_27;
  wire  _T_28;
  wire  _T_29;
  wire  RetimeWrapper_1_clock;
  wire  RetimeWrapper_1_reset;
  wire  RetimeWrapper_1_io_flow;
  wire  RetimeWrapper_1_io_in;
  wire  RetimeWrapper_1_io_out;
  wire  _T_33;
  wire  _T_34;
  wire  RetimeWrapper_2_clock;
  wire  RetimeWrapper_2_reset;
  wire  RetimeWrapper_2_io_flow;
  wire  RetimeWrapper_2_io_in;
  wire  RetimeWrapper_2_io_out;
  wire  _T_38;
  wire  RetimeWrapper_3_clock;
  wire  RetimeWrapper_3_reset;
  wire  RetimeWrapper_3_io_flow;
  wire  RetimeWrapper_3_io_in;
  wire  RetimeWrapper_3_io_out;
  wire  _T_42;
  wire  _T_43;
  wire  RetimeWrapper_4_clock;
  wire  RetimeWrapper_4_reset;
  wire  RetimeWrapper_4_io_flow;
  wire  RetimeWrapper_4_io_in;
  wire  RetimeWrapper_4_io_out;
  wire  _T_47;
  wire  _T_48;
  wire  _T_49;
  wire  _T_50;
  wire  _T_51;
  wire  RetimeWrapper_5_clock;
  wire  RetimeWrapper_5_reset;
  wire  RetimeWrapper_5_io_flow;
  wire  RetimeWrapper_5_io_in;
  wire  RetimeWrapper_5_io_out;
  wire  _T_55;
  wire  _T_56;
  wire  _T_57;
  wire  RetimeWrapper_6_clock;
  wire  RetimeWrapper_6_reset;
  wire  RetimeWrapper_6_io_flow;
  wire  RetimeWrapper_6_io_in;
  wire  RetimeWrapper_6_io_out;
  wire  _T_61;
  wire  _T_62;
  wire  RetimeWrapper_7_clock;
  wire  RetimeWrapper_7_reset;
  wire  RetimeWrapper_7_io_flow;
  wire  RetimeWrapper_7_io_in;
  wire  RetimeWrapper_7_io_out;
  wire  _T_66;
  wire  RetimeWrapper_8_clock;
  wire  RetimeWrapper_8_reset;
  wire  RetimeWrapper_8_io_flow;
  wire  RetimeWrapper_8_io_in;
  wire  RetimeWrapper_8_io_out;
  wire  _T_70;
  wire  _T_71;
  wire  RetimeWrapper_9_clock;
  wire  RetimeWrapper_9_reset;
  wire  RetimeWrapper_9_io_flow;
  wire  RetimeWrapper_9_io_in;
  wire  RetimeWrapper_9_io_out;
  wire  _T_75;
  wire  anyEnabled;
  wire  _T_76;
  wire  _T_77;
  wire  _T_78;
  wire  _T_79;
  wire  _T_80;
  wire  _T_81;
  wire  _T_82;
  reg  _T_85;
  reg [31:0] _RAND_0;
  wire  _T_91;
  wire  statesIn_0_clock;
  wire  statesIn_0_reset;
  wire  statesIn_0_io_input_enable;
  wire [1:0] statesIn_0_io_output_count;
  wire  statesOut_0_clock;
  wire  statesOut_0_reset;
  wire  statesOut_0_io_input_countUp;
  wire  statesOut_0_io_input_enable;
  wire [1:0] statesOut_0_io_output_count;
  wire  statesOut_1_clock;
  wire  statesOut_1_reset;
  wire  statesOut_1_io_input_countUp;
  wire  statesOut_1_io_input_enable;
  wire [1:0] statesOut_1_io_output_count;
  wire  _T_96;
  wire [31:0] _T_98_data;
  wire  _T_98_enable;
  wire  _T_98_reset;
  wire  _T_99;
  wire  _T_102;
  wire [31:0] _T_104_data;
  wire  _T_104_enable;
  wire  _T_104_reset;
  wire  _T_105;
  wire  _T_127;
  wire  _T_129;
  wire [31:0] _T_132_0;
  wire [31:0] _T_132_1;
  wire [31:0] _T_139;
  wire [31:0] _T_141;
  wire [31:0] _T_142;
  wire [31:0] _T_144;
  FF_1 ff_0 (
    .clock(ff_0_clock),
    .reset(ff_0_reset),
    .io_input_0_data(ff_0_io_input_0_data),
    .io_input_0_init(ff_0_io_input_0_init),
    .io_input_0_enable(ff_0_io_input_0_enable),
    .io_input_0_reset(ff_0_io_input_0_reset),
    .io_output_data(ff_0_io_output_data)
  );
  FF_1 ff_1 (
    .clock(ff_1_clock),
    .reset(ff_1_reset),
    .io_input_0_data(ff_1_io_input_0_data),
    .io_input_0_init(ff_1_io_input_0_init),
    .io_input_0_enable(ff_1_io_input_0_enable),
    .io_input_0_reset(ff_1_io_input_0_reset),
    .io_output_data(ff_1_io_output_data)
  );
  SRFF sEn_latch_0 (
    .clock(sEn_latch_0_clock),
    .reset(sEn_latch_0_reset),
    .io_input_set(sEn_latch_0_io_input_set),
    .io_input_reset(sEn_latch_0_io_input_reset),
    .io_input_asyn_reset(sEn_latch_0_io_input_asyn_reset),
    .io_output_data(sEn_latch_0_io_output_data)
  );
  SRFF sEn_latch_1 (
    .clock(sEn_latch_1_clock),
    .reset(sEn_latch_1_reset),
    .io_input_set(sEn_latch_1_io_input_set),
    .io_input_reset(sEn_latch_1_io_input_reset),
    .io_input_asyn_reset(sEn_latch_1_io_input_asyn_reset),
    .io_output_data(sEn_latch_1_io_output_data)
  );
  SRFF sDone_latch_0 (
    .clock(sDone_latch_0_clock),
    .reset(sDone_latch_0_reset),
    .io_input_set(sDone_latch_0_io_input_set),
    .io_input_reset(sDone_latch_0_io_input_reset),
    .io_input_asyn_reset(sDone_latch_0_io_input_asyn_reset),
    .io_output_data(sDone_latch_0_io_output_data)
  );
  SRFF sDone_latch_1 (
    .clock(sDone_latch_1_clock),
    .reset(sDone_latch_1_reset),
    .io_input_set(sDone_latch_1_io_input_set),
    .io_input_reset(sDone_latch_1_io_input_reset),
    .io_input_asyn_reset(sDone_latch_1_io_input_asyn_reset),
    .io_output_data(sDone_latch_1_io_output_data)
  );
  RetimeWrapper RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 (
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 (
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 (
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 (
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 (
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 (
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 (
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper RetimeWrapper_8 (
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper RetimeWrapper_9 (
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  NBufCtr_46 statesIn_0 (
    .clock(statesIn_0_clock),
    .reset(statesIn_0_reset),
    .io_input_enable(statesIn_0_io_input_enable),
    .io_output_count(statesIn_0_io_output_count)
  );
  NBufCtr_36 statesOut_0 (
    .clock(statesOut_0_clock),
    .reset(statesOut_0_reset),
    .io_input_countUp(statesOut_0_io_input_countUp),
    .io_input_enable(statesOut_0_io_input_enable),
    .io_output_count(statesOut_0_io_output_count)
  );
  NBufCtr_38 statesOut_1 (
    .clock(statesOut_1_clock),
    .reset(statesOut_1_reset),
    .io_input_countUp(statesOut_1_io_input_countUp),
    .io_input_enable(statesOut_1_io_input_enable),
    .io_output_count(statesOut_1_io_output_count)
  );
  assign _T_20 = ~ io_sDone_0;
  assign _T_21 = io_sEn_0 & _T_20;
  assign _T_22 = io_sEn_0 & io_sDone_0;
  assign _T_23 = ~ io_sEn_0;
  assign _T_28 = _T_22 & _T_27;
  assign _T_29 = _T_21 | _T_28;
  assign _T_34 = swap | _T_33;
  assign _T_43 = swap | _T_42;
  assign _T_48 = ~ io_sDone_1;
  assign _T_49 = io_sEn_1 & _T_48;
  assign _T_50 = io_sEn_1 & io_sDone_1;
  assign _T_51 = ~ io_sEn_1;
  assign _T_56 = _T_50 & _T_55;
  assign _T_57 = _T_49 | _T_56;
  assign _T_62 = swap | _T_61;
  assign _T_71 = swap | _T_70;
  assign anyEnabled = sEn_latch_0_io_output_data | sEn_latch_1_io_output_data;
  assign _T_76 = sDone_latch_0_io_output_data | io_sDone_0;
  assign _T_77 = sEn_latch_0_io_output_data == _T_76;
  assign _T_78 = sDone_latch_1_io_output_data | io_sDone_1;
  assign _T_79 = sEn_latch_1_io_output_data == _T_78;
  assign _T_80 = _T_77 & _T_79;
  assign _T_81 = _T_80 & anyEnabled;
  assign _T_82 = ~ _T_81;
  assign _T_91 = _T_81 & _T_85;
  assign _T_96 = statesIn_0_io_output_count == 2'h0;
  assign _T_99 = io_input_0_enable & _T_96;
  assign _T_102 = statesIn_0_io_output_count == 2'h1;
  assign _T_105 = io_input_0_enable & _T_102;
  assign _T_127 = statesOut_1_io_output_count == 2'h0;
  assign _T_129 = statesOut_1_io_output_count == 2'h1;
  assign _T_139 = _T_127 ? _T_132_0 : 32'h0;
  assign _T_141 = _T_129 ? _T_132_1 : 32'h0;
  assign _T_142 = _T_139 | _T_141;
  assign io_output_1_data = _T_144;
  assign ff_0_io_input_0_data = _T_98_data;
  assign ff_0_io_input_0_init = 32'h0;
  assign ff_0_io_input_0_enable = _T_98_enable;
  assign ff_0_io_input_0_reset = _T_98_reset;
  assign ff_0_clock = clock;
  assign ff_0_reset = reset;
  assign ff_1_io_input_0_data = _T_104_data;
  assign ff_1_io_input_0_init = 32'h0;
  assign ff_1_io_input_0_enable = _T_104_enable;
  assign ff_1_io_input_0_reset = _T_104_reset;
  assign ff_1_clock = clock;
  assign ff_1_reset = reset;
  assign sEn_latch_0_io_input_set = _T_29;
  assign sEn_latch_0_io_input_reset = _T_34;
  assign sEn_latch_0_io_input_asyn_reset = _T_38;
  assign sEn_latch_0_clock = clock;
  assign sEn_latch_0_reset = reset;
  assign sEn_latch_1_io_input_set = _T_57;
  assign sEn_latch_1_io_input_reset = _T_62;
  assign sEn_latch_1_io_input_asyn_reset = _T_66;
  assign sEn_latch_1_clock = clock;
  assign sEn_latch_1_reset = reset;
  assign sDone_latch_0_io_input_set = io_sDone_0;
  assign sDone_latch_0_io_input_reset = _T_43;
  assign sDone_latch_0_io_input_asyn_reset = _T_47;
  assign sDone_latch_0_clock = clock;
  assign sDone_latch_0_reset = reset;
  assign sDone_latch_1_io_input_set = io_sDone_1;
  assign sDone_latch_1_io_input_reset = _T_71;
  assign sDone_latch_1_io_input_asyn_reset = _T_75;
  assign sDone_latch_1_clock = clock;
  assign sDone_latch_1_reset = reset;
  assign swap = _T_91;
  assign RetimeWrapper_io_flow = 1'h1;
  assign RetimeWrapper_io_in = _T_23;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_27 = RetimeWrapper_io_out;
  assign RetimeWrapper_1_io_flow = 1'h1;
  assign RetimeWrapper_1_io_in = swap;
  assign RetimeWrapper_1_clock = clock;
  assign RetimeWrapper_1_reset = reset;
  assign _T_33 = RetimeWrapper_1_io_out;
  assign RetimeWrapper_2_io_flow = 1'h1;
  assign RetimeWrapper_2_io_in = reset;
  assign RetimeWrapper_2_clock = clock;
  assign RetimeWrapper_2_reset = reset;
  assign _T_38 = RetimeWrapper_2_io_out;
  assign RetimeWrapper_3_io_flow = 1'h1;
  assign RetimeWrapper_3_io_in = swap;
  assign RetimeWrapper_3_clock = clock;
  assign RetimeWrapper_3_reset = reset;
  assign _T_42 = RetimeWrapper_3_io_out;
  assign RetimeWrapper_4_io_flow = 1'h1;
  assign RetimeWrapper_4_io_in = reset;
  assign RetimeWrapper_4_clock = clock;
  assign RetimeWrapper_4_reset = reset;
  assign _T_47 = RetimeWrapper_4_io_out;
  assign RetimeWrapper_5_io_flow = 1'h1;
  assign RetimeWrapper_5_io_in = _T_51;
  assign RetimeWrapper_5_clock = clock;
  assign RetimeWrapper_5_reset = reset;
  assign _T_55 = RetimeWrapper_5_io_out;
  assign RetimeWrapper_6_io_flow = 1'h1;
  assign RetimeWrapper_6_io_in = swap;
  assign RetimeWrapper_6_clock = clock;
  assign RetimeWrapper_6_reset = reset;
  assign _T_61 = RetimeWrapper_6_io_out;
  assign RetimeWrapper_7_io_flow = 1'h1;
  assign RetimeWrapper_7_io_in = reset;
  assign RetimeWrapper_7_clock = clock;
  assign RetimeWrapper_7_reset = reset;
  assign _T_66 = RetimeWrapper_7_io_out;
  assign RetimeWrapper_8_io_flow = 1'h1;
  assign RetimeWrapper_8_io_in = swap;
  assign RetimeWrapper_8_clock = clock;
  assign RetimeWrapper_8_reset = reset;
  assign _T_70 = RetimeWrapper_8_io_out;
  assign RetimeWrapper_9_io_flow = 1'h1;
  assign RetimeWrapper_9_io_in = reset;
  assign RetimeWrapper_9_clock = clock;
  assign RetimeWrapper_9_reset = reset;
  assign _T_75 = RetimeWrapper_9_io_out;
  assign statesIn_0_io_input_enable = swap;
  assign statesIn_0_clock = clock;
  assign statesIn_0_reset = reset;
  assign statesOut_0_io_input_countUp = 1'h0;
  assign statesOut_0_io_input_enable = swap;
  assign statesOut_0_clock = clock;
  assign statesOut_0_reset = reset;
  assign statesOut_1_io_input_countUp = 1'h0;
  assign statesOut_1_io_input_enable = swap;
  assign statesOut_1_clock = clock;
  assign statesOut_1_reset = reset;
  assign _T_98_data = io_input_0_data;
  assign _T_98_enable = _T_99;
  assign _T_98_reset = io_input_0_reset;
  assign _T_104_data = io_input_0_data;
  assign _T_104_enable = _T_105;
  assign _T_104_reset = io_input_0_reset;
  assign _T_132_0 = ff_0_io_output_data;
  assign _T_132_1 = ff_1_io_output_data;
  assign _T_144 = _T_142;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_85 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_85 <= 1'h0;
    end else begin
      _T_85 <= _T_82;
    end
  end
endmodule
module SingleCounter_17(
  input         clock,
  input         reset,
  input  [31:0] io_input_stop,
  input         io_input_reset,
  input         io_input_enable,
  output [31:0] io_output_count_0,
  output [31:0] io_output_count_1,
  output [31:0] io_output_count_2,
  output [31:0] io_output_count_3,
  output        io_output_done
);
  wire  FF_clock;
  wire  FF_reset;
  wire [31:0] FF_io_input_0_data;
  wire [31:0] FF_io_input_0_init;
  wire  FF_io_input_0_enable;
  wire  FF_io_input_0_reset;
  wire [31:0] FF_io_output_data;
  wire  FF_1_clock;
  wire  FF_1_reset;
  wire [31:0] FF_1_io_input_0_data;
  wire [31:0] FF_1_io_input_0_init;
  wire  FF_1_io_input_0_enable;
  wire  FF_1_io_input_0_reset;
  wire [31:0] FF_1_io_output_data;
  wire  FF_2_clock;
  wire  FF_2_reset;
  wire [31:0] FF_2_io_input_0_data;
  wire [31:0] FF_2_io_input_0_init;
  wire  FF_2_io_input_0_enable;
  wire  FF_2_io_input_0_reset;
  wire [31:0] FF_2_io_output_data;
  wire  FF_3_clock;
  wire  FF_3_reset;
  wire [31:0] FF_3_io_input_0_data;
  wire [31:0] FF_3_io_input_0_init;
  wire  FF_3_io_input_0_enable;
  wire  FF_3_io_input_0_reset;
  wire [31:0] FF_3_io_output_data;
  wire [31:0] _T_30;
  wire [31:0] _T_31;
  wire [31:0] _T_32;
  wire [31:0] _T_33;
  wire [32:0] _T_35;
  wire [31:0] _T_36;
  wire [31:0] _T_37;
  wire [32:0] _T_38;
  wire [31:0] _T_39;
  wire [31:0] _T_40;
  wire [32:0] _T_41;
  wire [31:0] _T_42;
  wire [31:0] _T_43;
  wire [32:0] _T_44;
  wire [31:0] _T_45;
  wire [31:0] _T_46;
  wire  _T_49;
  wire [31:0] _T_62;
  wire [31:0] _T_63;
  wire [31:0] _T_64;
  wire [31:0] _T_69;
  wire [31:0] _T_70;
  wire [31:0] _T_71;
  wire [31:0] _T_76;
  wire [31:0] _T_77;
  wire [31:0] _T_78;
  wire [31:0] _T_83;
  wire [31:0] _T_84;
  wire [31:0] _T_85;
  wire  _T_98;
  FF_1 FF (
    .clock(FF_clock),
    .reset(FF_reset),
    .io_input_0_data(FF_io_input_0_data),
    .io_input_0_init(FF_io_input_0_init),
    .io_input_0_enable(FF_io_input_0_enable),
    .io_input_0_reset(FF_io_input_0_reset),
    .io_output_data(FF_io_output_data)
  );
  FF_1 FF_1 (
    .clock(FF_1_clock),
    .reset(FF_1_reset),
    .io_input_0_data(FF_1_io_input_0_data),
    .io_input_0_init(FF_1_io_input_0_init),
    .io_input_0_enable(FF_1_io_input_0_enable),
    .io_input_0_reset(FF_1_io_input_0_reset),
    .io_output_data(FF_1_io_output_data)
  );
  FF_1 FF_2 (
    .clock(FF_2_clock),
    .reset(FF_2_reset),
    .io_input_0_data(FF_2_io_input_0_data),
    .io_input_0_init(FF_2_io_input_0_init),
    .io_input_0_enable(FF_2_io_input_0_enable),
    .io_input_0_reset(FF_2_io_input_0_reset),
    .io_output_data(FF_2_io_output_data)
  );
  FF_1 FF_3 (
    .clock(FF_3_clock),
    .reset(FF_3_reset),
    .io_input_0_data(FF_3_io_input_0_data),
    .io_input_0_init(FF_3_io_input_0_init),
    .io_input_0_enable(FF_3_io_input_0_enable),
    .io_input_0_reset(FF_3_io_input_0_reset),
    .io_output_data(FF_3_io_output_data)
  );
  assign _T_30 = $signed(FF_io_output_data);
  assign _T_31 = $signed(FF_1_io_output_data);
  assign _T_32 = $signed(FF_2_io_output_data);
  assign _T_33 = $signed(FF_3_io_output_data);
  assign _T_35 = $signed(_T_30) + $signed(32'sh4);
  assign _T_36 = _T_35[31:0];
  assign _T_37 = $signed(_T_36);
  assign _T_38 = $signed(_T_31) + $signed(32'sh4);
  assign _T_39 = _T_38[31:0];
  assign _T_40 = $signed(_T_39);
  assign _T_41 = $signed(_T_32) + $signed(32'sh4);
  assign _T_42 = _T_41[31:0];
  assign _T_43 = $signed(_T_42);
  assign _T_44 = $signed(_T_33) + $signed(32'sh4);
  assign _T_45 = _T_44[31:0];
  assign _T_46 = $signed(_T_45);
  assign _T_49 = $signed(_T_37) >= $signed(io_input_stop);
  assign _T_62 = $unsigned(_T_37);
  assign _T_63 = _T_49 ? 32'h0 : _T_62;
  assign _T_64 = io_input_reset ? 32'h0 : _T_63;
  assign _T_69 = $unsigned(_T_40);
  assign _T_70 = _T_49 ? 32'h1 : _T_69;
  assign _T_71 = io_input_reset ? 32'h1 : _T_70;
  assign _T_76 = $unsigned(_T_43);
  assign _T_77 = _T_49 ? 32'h2 : _T_76;
  assign _T_78 = io_input_reset ? 32'h2 : _T_77;
  assign _T_83 = $unsigned(_T_46);
  assign _T_84 = _T_49 ? 32'h3 : _T_83;
  assign _T_85 = io_input_reset ? 32'h3 : _T_84;
  assign _T_98 = io_input_enable & _T_49;
  assign io_output_count_0 = _T_30;
  assign io_output_count_1 = _T_31;
  assign io_output_count_2 = _T_32;
  assign io_output_count_3 = _T_33;
  assign io_output_done = _T_98;
  assign FF_io_input_0_data = _T_64;
  assign FF_io_input_0_init = 32'h0;
  assign FF_io_input_0_enable = io_input_enable;
  assign FF_io_input_0_reset = io_input_reset;
  assign FF_clock = clock;
  assign FF_reset = reset;
  assign FF_1_io_input_0_data = _T_71;
  assign FF_1_io_input_0_init = 32'h1;
  assign FF_1_io_input_0_enable = io_input_enable;
  assign FF_1_io_input_0_reset = io_input_reset;
  assign FF_1_clock = clock;
  assign FF_1_reset = reset;
  assign FF_2_io_input_0_data = _T_78;
  assign FF_2_io_input_0_init = 32'h2;
  assign FF_2_io_input_0_enable = io_input_enable;
  assign FF_2_io_input_0_reset = io_input_reset;
  assign FF_2_clock = clock;
  assign FF_2_reset = reset;
  assign FF_3_io_input_0_data = _T_85;
  assign FF_3_io_input_0_init = 32'h3;
  assign FF_3_io_input_0_enable = io_input_enable;
  assign FF_3_io_input_0_reset = io_input_reset;
  assign FF_3_clock = clock;
  assign FF_3_reset = reset;
endmodule
module Counter_5(
  input         clock,
  input         reset,
  input  [31:0] io_input_stops_0,
  input         io_input_reset,
  input         io_input_enable,
  output [31:0] io_output_counts_3,
  output [31:0] io_output_counts_2,
  output [31:0] io_output_counts_1,
  output [31:0] io_output_counts_0,
  output        io_output_done
);
  wire  ctrs_0_clock;
  wire  ctrs_0_reset;
  wire [31:0] ctrs_0_io_input_stop;
  wire  ctrs_0_io_input_reset;
  wire  ctrs_0_io_input_enable;
  wire [31:0] ctrs_0_io_output_count_0;
  wire [31:0] ctrs_0_io_output_count_1;
  wire [31:0] ctrs_0_io_output_count_2;
  wire [31:0] ctrs_0_io_output_count_3;
  wire  ctrs_0_io_output_done;
  reg  wasDone;
  reg [31:0] _RAND_0;
  wire  _T_35;
  wire  _T_36;
  wire  _T_37;
  SingleCounter_17 ctrs_0 (
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_input_stop(ctrs_0_io_input_stop),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_count_1(ctrs_0_io_output_count_1),
    .io_output_count_2(ctrs_0_io_output_count_2),
    .io_output_count_3(ctrs_0_io_output_count_3),
    .io_output_done(ctrs_0_io_output_done)
  );
  assign _T_35 = io_input_enable & ctrs_0_io_output_done;
  assign _T_36 = ~ wasDone;
  assign _T_37 = _T_35 & _T_36;
  assign io_output_counts_3 = ctrs_0_io_output_count_3;
  assign io_output_counts_2 = ctrs_0_io_output_count_2;
  assign io_output_counts_1 = ctrs_0_io_output_count_1;
  assign io_output_counts_0 = ctrs_0_io_output_count_0;
  assign io_output_done = _T_37;
  assign ctrs_0_io_input_stop = io_input_stops_0;
  assign ctrs_0_io_input_reset = io_input_reset;
  assign ctrs_0_io_input_enable = io_input_enable;
  assign ctrs_0_clock = clock;
  assign ctrs_0_reset = reset;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= ctrs_0_io_output_done;
    end
  end
endmodule
module Innerpipe_10(
  input   clock,
  input   reset,
  input   io_input_enable,
  input   io_input_ctr_done,
  input   io_input_rst,
  output  io_output_done,
  output  io_output_ctr_inc,
  output  io_output_rst_en
);
  wire  SRFF_clock;
  wire  SRFF_reset;
  wire  SRFF_io_input_set;
  wire  SRFF_io_input_reset;
  wire  SRFF_io_input_asyn_reset;
  wire  SRFF_io_output_data;
  wire  FF_clock;
  wire  FF_reset;
  wire [31:0] FF_io_input_0_data;
  wire [31:0] FF_io_input_0_init;
  wire  FF_io_input_0_enable;
  wire  FF_io_input_0_reset;
  wire [31:0] FF_io_output_data;
  wire  _T_19;
  wire  _T_20;
  wire  _T_22;
  wire  _T_24;
  wire  _T_25;
  wire  _T_26;
  wire  _T_28;
  wire  _T_31;
  wire  _T_32;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire  RetimeWrapper_io_flow;
  wire  RetimeWrapper_io_in;
  wire  RetimeWrapper_io_out;
  wire  _T_36;
  wire  _T_37;
  wire  _T_39;
  wire [1:0] _T_45;
  wire [1:0] _T_48;
  wire [1:0] _GEN_0;
  wire  _T_50;
  wire  _T_53;
  wire  RetimeWrapper_1_clock;
  wire  RetimeWrapper_1_reset;
  wire  RetimeWrapper_1_io_flow;
  wire  RetimeWrapper_1_io_in;
  wire  RetimeWrapper_1_io_out;
  wire  _T_57;
  wire  _T_58;
  wire  _T_59;
  wire  _T_60;
  wire  _GEN_3;
  wire  _T_76;
  wire  _T_84;
  wire [32:0] _T_92;
  wire [31:0] _T_93;
  wire [31:0] _T_94;
  wire [31:0] _GEN_9;
  wire  _GEN_10;
  wire  _GEN_11;
  wire [31:0] _GEN_13;
  wire  _GEN_14;
  wire  _GEN_16;
  wire [31:0] _GEN_17;
  wire  _T_97;
  wire  _T_98;
  wire  _GEN_18;
  wire  _GEN_20;
  wire [31:0] _GEN_21;
  SRFF SRFF (
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output_data(SRFF_io_output_data)
  );
  FF_1 FF (
    .clock(FF_clock),
    .reset(FF_reset),
    .io_input_0_data(FF_io_input_0_data),
    .io_input_0_init(FF_io_input_0_init),
    .io_input_0_enable(FF_io_input_0_enable),
    .io_input_0_reset(FF_io_input_0_reset),
    .io_output_data(FF_io_output_data)
  );
  RetimeWrapper RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 (
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign _T_19 = ~ io_input_enable;
  assign _T_20 = _T_19 | io_input_rst;
  assign _T_22 = FF_io_output_data != 32'h3;
  assign _T_24 = FF_io_output_data != 32'h1;
  assign _T_25 = _T_22 & _T_24;
  assign _T_26 = _T_20 | _T_25;
  assign _T_28 = FF_io_output_data != 32'h2;
  assign _T_31 = _T_28 & _T_24;
  assign _T_32 = _T_31 | SRFF_io_output_data;
  assign _T_37 = _T_36 | io_input_rst;
  assign _T_39 = FF_io_output_data == 32'h1;
  assign _T_45 = io_input_ctr_done ? 2'h3 : 2'h2;
  assign _T_48 = io_input_ctr_done ? 2'h3 : 2'h1;
  assign _GEN_0 = _T_26 ? _T_48 : _T_45;
  assign _T_50 = FF_io_output_data == 32'h2;
  assign _T_53 = _T_28 | SRFF_io_output_data;
  assign _T_58 = _T_57 | io_input_rst;
  assign _T_59 = ~ _T_58;
  assign _T_60 = io_input_enable & _T_59;
  assign _GEN_3 = io_input_ctr_done ? 1'h0 : _T_60;
  assign _T_76 = FF_io_output_data == 32'h3;
  assign _T_84 = FF_io_output_data >= 32'h4;
  assign _T_92 = FF_io_output_data + 32'h1;
  assign _T_93 = _T_92[31:0];
  assign _T_94 = _T_84 ? 32'h1 : _T_93;
  assign _GEN_9 = _T_76 ? 32'h1 : _T_94;
  assign _GEN_10 = _T_50 ? _GEN_3 : 1'h0;
  assign _GEN_11 = _T_50 ? io_input_ctr_done : 1'h0;
  assign _GEN_13 = _T_50 ? {{30'd0}, _T_45} : _GEN_9;
  assign _GEN_14 = _T_39 ? 1'h0 : _GEN_11;
  assign _GEN_16 = _T_39 ? 1'h0 : _GEN_10;
  assign _GEN_17 = _T_39 ? {{30'd0}, _GEN_0} : _GEN_13;
  assign _T_97 = _T_50 & io_input_ctr_done;
  assign _T_98 = io_input_ctr_done | _T_97;
  assign _GEN_18 = io_input_enable ? _GEN_14 : _T_98;
  assign _GEN_20 = io_input_enable ? _GEN_16 : 1'h0;
  assign _GEN_21 = io_input_enable ? _GEN_17 : 32'h1;
  assign io_output_done = _GEN_18;
  assign io_output_ctr_inc = _GEN_20;
  assign io_output_rst_en = _T_37;
  assign SRFF_io_input_set = io_input_rst;
  assign SRFF_io_input_reset = io_input_enable;
  assign SRFF_io_input_asyn_reset = io_input_enable;
  assign SRFF_clock = clock;
  assign SRFF_reset = reset;
  assign FF_io_input_0_data = _GEN_21;
  assign FF_io_input_0_init = 32'h1;
  assign FF_io_input_0_enable = 1'h1;
  assign FF_io_input_0_reset = 1'h0;
  assign FF_clock = clock;
  assign FF_reset = reset;
  assign RetimeWrapper_io_flow = 1'h1;
  assign RetimeWrapper_io_in = _T_32;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_36 = RetimeWrapper_io_out;
  assign RetimeWrapper_1_io_flow = 1'h1;
  assign RetimeWrapper_1_io_in = _T_53;
  assign RetimeWrapper_1_clock = clock;
  assign RetimeWrapper_1_reset = reset;
  assign _T_57 = RetimeWrapper_1_io_out;
endmodule
module FF_103(
  input   clock,
  input   reset,
  input   io_input_0_data,
  input   io_input_0_enable,
  input   io_input_0_reset,
  output  io_output_data
);
  reg  ff;
  reg [31:0] _RAND_0;
  wire  _T_7;
  wire  _T_8;
  wire  _T_9;
  assign _T_7 = io_input_0_enable ? io_input_0_data : ff;
  assign _T_8 = io_input_0_reset ? 1'h0 : _T_7;
  assign _T_9 = io_input_0_reset ? 1'h0 : ff;
  assign io_output_data = _T_9;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  ff = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 1'h0;
    end else begin
      if (io_input_0_reset) begin
        ff <= 1'h0;
      end else begin
        if (io_input_0_enable) begin
          ff <= io_input_0_data;
        end
      end
    end
  end
endmodule
module NBufFF_6(
  input   clock,
  input   reset,
  input   io_sEn_0,
  input   io_sEn_1,
  input   io_sEn_2,
  input   io_sEn_3,
  input   io_sEn_4,
  input   io_sDone_0,
  input   io_sDone_1,
  input   io_sDone_2,
  input   io_sDone_3,
  input   io_sDone_4,
  input   io_input_0_data,
  input   io_input_0_enable,
  input   io_input_0_reset,
  output  io_output_1_data,
  output  io_output_2_data,
  output  io_output_3_data,
  output  io_output_4_data
);
  wire  ff_0_clock;
  wire  ff_0_reset;
  wire  ff_0_io_input_0_data;
  wire  ff_0_io_input_0_enable;
  wire  ff_0_io_input_0_reset;
  wire  ff_0_io_output_data;
  wire  ff_1_clock;
  wire  ff_1_reset;
  wire  ff_1_io_input_0_data;
  wire  ff_1_io_input_0_enable;
  wire  ff_1_io_input_0_reset;
  wire  ff_1_io_output_data;
  wire  ff_2_clock;
  wire  ff_2_reset;
  wire  ff_2_io_input_0_data;
  wire  ff_2_io_input_0_enable;
  wire  ff_2_io_input_0_reset;
  wire  ff_2_io_output_data;
  wire  ff_3_clock;
  wire  ff_3_reset;
  wire  ff_3_io_input_0_data;
  wire  ff_3_io_input_0_enable;
  wire  ff_3_io_input_0_reset;
  wire  ff_3_io_output_data;
  wire  ff_4_clock;
  wire  ff_4_reset;
  wire  ff_4_io_input_0_data;
  wire  ff_4_io_input_0_enable;
  wire  ff_4_io_input_0_reset;
  wire  ff_4_io_output_data;
  wire  sEn_latch_0_clock;
  wire  sEn_latch_0_reset;
  wire  sEn_latch_0_io_input_set;
  wire  sEn_latch_0_io_input_reset;
  wire  sEn_latch_0_io_input_asyn_reset;
  wire  sEn_latch_0_io_output_data;
  wire  sEn_latch_1_clock;
  wire  sEn_latch_1_reset;
  wire  sEn_latch_1_io_input_set;
  wire  sEn_latch_1_io_input_reset;
  wire  sEn_latch_1_io_input_asyn_reset;
  wire  sEn_latch_1_io_output_data;
  wire  sEn_latch_2_clock;
  wire  sEn_latch_2_reset;
  wire  sEn_latch_2_io_input_set;
  wire  sEn_latch_2_io_input_reset;
  wire  sEn_latch_2_io_input_asyn_reset;
  wire  sEn_latch_2_io_output_data;
  wire  sEn_latch_3_clock;
  wire  sEn_latch_3_reset;
  wire  sEn_latch_3_io_input_set;
  wire  sEn_latch_3_io_input_reset;
  wire  sEn_latch_3_io_input_asyn_reset;
  wire  sEn_latch_3_io_output_data;
  wire  sEn_latch_4_clock;
  wire  sEn_latch_4_reset;
  wire  sEn_latch_4_io_input_set;
  wire  sEn_latch_4_io_input_reset;
  wire  sEn_latch_4_io_input_asyn_reset;
  wire  sEn_latch_4_io_output_data;
  wire  sDone_latch_0_clock;
  wire  sDone_latch_0_reset;
  wire  sDone_latch_0_io_input_set;
  wire  sDone_latch_0_io_input_reset;
  wire  sDone_latch_0_io_input_asyn_reset;
  wire  sDone_latch_0_io_output_data;
  wire  sDone_latch_1_clock;
  wire  sDone_latch_1_reset;
  wire  sDone_latch_1_io_input_set;
  wire  sDone_latch_1_io_input_reset;
  wire  sDone_latch_1_io_input_asyn_reset;
  wire  sDone_latch_1_io_output_data;
  wire  sDone_latch_2_clock;
  wire  sDone_latch_2_reset;
  wire  sDone_latch_2_io_input_set;
  wire  sDone_latch_2_io_input_reset;
  wire  sDone_latch_2_io_input_asyn_reset;
  wire  sDone_latch_2_io_output_data;
  wire  sDone_latch_3_clock;
  wire  sDone_latch_3_reset;
  wire  sDone_latch_3_io_input_set;
  wire  sDone_latch_3_io_input_reset;
  wire  sDone_latch_3_io_input_asyn_reset;
  wire  sDone_latch_3_io_output_data;
  wire  sDone_latch_4_clock;
  wire  sDone_latch_4_reset;
  wire  sDone_latch_4_io_input_set;
  wire  sDone_latch_4_io_input_reset;
  wire  sDone_latch_4_io_input_asyn_reset;
  wire  sDone_latch_4_io_output_data;
  wire  swap;
  wire  _T_20;
  wire  _T_21;
  wire  _T_22;
  wire  _T_23;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire  RetimeWrapper_io_flow;
  wire  RetimeWrapper_io_in;
  wire  RetimeWrapper_io_out;
  wire  _T_27;
  wire  _T_28;
  wire  _T_29;
  wire  RetimeWrapper_1_clock;
  wire  RetimeWrapper_1_reset;
  wire  RetimeWrapper_1_io_flow;
  wire  RetimeWrapper_1_io_in;
  wire  RetimeWrapper_1_io_out;
  wire  _T_33;
  wire  _T_34;
  wire  RetimeWrapper_2_clock;
  wire  RetimeWrapper_2_reset;
  wire  RetimeWrapper_2_io_flow;
  wire  RetimeWrapper_2_io_in;
  wire  RetimeWrapper_2_io_out;
  wire  _T_38;
  wire  RetimeWrapper_3_clock;
  wire  RetimeWrapper_3_reset;
  wire  RetimeWrapper_3_io_flow;
  wire  RetimeWrapper_3_io_in;
  wire  RetimeWrapper_3_io_out;
  wire  _T_42;
  wire  _T_43;
  wire  RetimeWrapper_4_clock;
  wire  RetimeWrapper_4_reset;
  wire  RetimeWrapper_4_io_flow;
  wire  RetimeWrapper_4_io_in;
  wire  RetimeWrapper_4_io_out;
  wire  _T_47;
  wire  _T_48;
  wire  _T_49;
  wire  _T_50;
  wire  _T_51;
  wire  RetimeWrapper_5_clock;
  wire  RetimeWrapper_5_reset;
  wire  RetimeWrapper_5_io_flow;
  wire  RetimeWrapper_5_io_in;
  wire  RetimeWrapper_5_io_out;
  wire  _T_55;
  wire  _T_56;
  wire  _T_57;
  wire  RetimeWrapper_6_clock;
  wire  RetimeWrapper_6_reset;
  wire  RetimeWrapper_6_io_flow;
  wire  RetimeWrapper_6_io_in;
  wire  RetimeWrapper_6_io_out;
  wire  _T_61;
  wire  _T_62;
  wire  RetimeWrapper_7_clock;
  wire  RetimeWrapper_7_reset;
  wire  RetimeWrapper_7_io_flow;
  wire  RetimeWrapper_7_io_in;
  wire  RetimeWrapper_7_io_out;
  wire  _T_66;
  wire  RetimeWrapper_8_clock;
  wire  RetimeWrapper_8_reset;
  wire  RetimeWrapper_8_io_flow;
  wire  RetimeWrapper_8_io_in;
  wire  RetimeWrapper_8_io_out;
  wire  _T_70;
  wire  _T_71;
  wire  RetimeWrapper_9_clock;
  wire  RetimeWrapper_9_reset;
  wire  RetimeWrapper_9_io_flow;
  wire  RetimeWrapper_9_io_in;
  wire  RetimeWrapper_9_io_out;
  wire  _T_75;
  wire  _T_76;
  wire  _T_77;
  wire  _T_78;
  wire  _T_79;
  wire  RetimeWrapper_10_clock;
  wire  RetimeWrapper_10_reset;
  wire  RetimeWrapper_10_io_flow;
  wire  RetimeWrapper_10_io_in;
  wire  RetimeWrapper_10_io_out;
  wire  _T_83;
  wire  _T_84;
  wire  _T_85;
  wire  RetimeWrapper_11_clock;
  wire  RetimeWrapper_11_reset;
  wire  RetimeWrapper_11_io_flow;
  wire  RetimeWrapper_11_io_in;
  wire  RetimeWrapper_11_io_out;
  wire  _T_89;
  wire  _T_90;
  wire  RetimeWrapper_12_clock;
  wire  RetimeWrapper_12_reset;
  wire  RetimeWrapper_12_io_flow;
  wire  RetimeWrapper_12_io_in;
  wire  RetimeWrapper_12_io_out;
  wire  _T_94;
  wire  RetimeWrapper_13_clock;
  wire  RetimeWrapper_13_reset;
  wire  RetimeWrapper_13_io_flow;
  wire  RetimeWrapper_13_io_in;
  wire  RetimeWrapper_13_io_out;
  wire  _T_98;
  wire  _T_99;
  wire  RetimeWrapper_14_clock;
  wire  RetimeWrapper_14_reset;
  wire  RetimeWrapper_14_io_flow;
  wire  RetimeWrapper_14_io_in;
  wire  RetimeWrapper_14_io_out;
  wire  _T_103;
  wire  _T_104;
  wire  _T_105;
  wire  _T_106;
  wire  _T_107;
  wire  RetimeWrapper_15_clock;
  wire  RetimeWrapper_15_reset;
  wire  RetimeWrapper_15_io_flow;
  wire  RetimeWrapper_15_io_in;
  wire  RetimeWrapper_15_io_out;
  wire  _T_111;
  wire  _T_112;
  wire  _T_113;
  wire  RetimeWrapper_16_clock;
  wire  RetimeWrapper_16_reset;
  wire  RetimeWrapper_16_io_flow;
  wire  RetimeWrapper_16_io_in;
  wire  RetimeWrapper_16_io_out;
  wire  _T_117;
  wire  _T_118;
  wire  RetimeWrapper_17_clock;
  wire  RetimeWrapper_17_reset;
  wire  RetimeWrapper_17_io_flow;
  wire  RetimeWrapper_17_io_in;
  wire  RetimeWrapper_17_io_out;
  wire  _T_122;
  wire  RetimeWrapper_18_clock;
  wire  RetimeWrapper_18_reset;
  wire  RetimeWrapper_18_io_flow;
  wire  RetimeWrapper_18_io_in;
  wire  RetimeWrapper_18_io_out;
  wire  _T_126;
  wire  _T_127;
  wire  RetimeWrapper_19_clock;
  wire  RetimeWrapper_19_reset;
  wire  RetimeWrapper_19_io_flow;
  wire  RetimeWrapper_19_io_in;
  wire  RetimeWrapper_19_io_out;
  wire  _T_131;
  wire  _T_132;
  wire  _T_133;
  wire  _T_134;
  wire  _T_135;
  wire  RetimeWrapper_20_clock;
  wire  RetimeWrapper_20_reset;
  wire  RetimeWrapper_20_io_flow;
  wire  RetimeWrapper_20_io_in;
  wire  RetimeWrapper_20_io_out;
  wire  _T_139;
  wire  _T_140;
  wire  _T_141;
  wire  RetimeWrapper_21_clock;
  wire  RetimeWrapper_21_reset;
  wire  RetimeWrapper_21_io_flow;
  wire  RetimeWrapper_21_io_in;
  wire  RetimeWrapper_21_io_out;
  wire  _T_145;
  wire  _T_146;
  wire  RetimeWrapper_22_clock;
  wire  RetimeWrapper_22_reset;
  wire  RetimeWrapper_22_io_flow;
  wire  RetimeWrapper_22_io_in;
  wire  RetimeWrapper_22_io_out;
  wire  _T_150;
  wire  RetimeWrapper_23_clock;
  wire  RetimeWrapper_23_reset;
  wire  RetimeWrapper_23_io_flow;
  wire  RetimeWrapper_23_io_in;
  wire  RetimeWrapper_23_io_out;
  wire  _T_154;
  wire  _T_155;
  wire  RetimeWrapper_24_clock;
  wire  RetimeWrapper_24_reset;
  wire  RetimeWrapper_24_io_flow;
  wire  RetimeWrapper_24_io_in;
  wire  RetimeWrapper_24_io_out;
  wire  _T_159;
  wire  _T_160;
  wire  _T_161;
  wire  _T_162;
  wire  anyEnabled;
  wire  _T_163;
  wire  _T_164;
  wire  _T_165;
  wire  _T_166;
  wire  _T_167;
  wire  _T_168;
  wire  _T_169;
  wire  _T_170;
  wire  _T_171;
  wire  _T_172;
  wire  _T_173;
  wire  _T_174;
  wire  _T_175;
  wire  _T_176;
  wire  _T_177;
  wire  _T_178;
  reg  _T_181;
  reg [31:0] _RAND_0;
  wire  _T_187;
  wire  statesIn_0_clock;
  wire  statesIn_0_reset;
  wire  statesIn_0_io_input_enable;
  wire [3:0] statesIn_0_io_output_count;
  wire  statesOut_0_clock;
  wire  statesOut_0_reset;
  wire  statesOut_0_io_input_enable;
  wire  statesOut_1_clock;
  wire  statesOut_1_reset;
  wire  statesOut_1_io_input_enable;
  wire [3:0] statesOut_1_io_output_count;
  wire  statesOut_2_clock;
  wire  statesOut_2_reset;
  wire  statesOut_2_io_input_enable;
  wire [3:0] statesOut_2_io_output_count;
  wire  statesOut_3_clock;
  wire  statesOut_3_reset;
  wire  statesOut_3_io_input_enable;
  wire [3:0] statesOut_3_io_output_count;
  wire  statesOut_4_clock;
  wire  statesOut_4_reset;
  wire  statesOut_4_io_input_enable;
  wire [3:0] statesOut_4_io_output_count;
  wire  _T_195;
  wire  _T_197_data;
  wire  _T_197_enable;
  wire  _T_197_reset;
  wire  _T_198;
  wire  _T_201;
  wire  _T_203_data;
  wire  _T_203_enable;
  wire  _T_203_reset;
  wire  _T_204;
  wire  _T_207;
  wire  _T_209_data;
  wire  _T_209_enable;
  wire  _T_209_reset;
  wire  _T_210;
  wire  _T_213;
  wire  _T_215_data;
  wire  _T_215_enable;
  wire  _T_215_reset;
  wire  _T_216;
  wire  _T_219;
  wire  _T_221_data;
  wire  _T_221_enable;
  wire  _T_221_reset;
  wire  _T_222;
  wire  _T_262;
  wire  _T_264;
  wire  _T_266;
  wire  _T_268;
  wire  _T_270;
  wire  _T_273_0;
  wire  _T_273_1;
  wire  _T_273_2;
  wire  _T_273_3;
  wire  _T_273_4;
  wire  _T_283;
  wire  _T_285;
  wire  _T_287;
  wire  _T_289;
  wire  _T_291;
  wire  _T_292;
  wire  _T_293;
  wire  _T_294;
  wire  _T_295;
  wire  _T_297;
  wire  _T_299;
  wire  _T_301;
  wire  _T_303;
  wire  _T_305;
  wire  _T_307;
  wire  _T_310_0;
  wire  _T_310_1;
  wire  _T_310_2;
  wire  _T_310_3;
  wire  _T_310_4;
  wire  _T_320;
  wire  _T_322;
  wire  _T_324;
  wire  _T_326;
  wire  _T_328;
  wire  _T_329;
  wire  _T_330;
  wire  _T_331;
  wire  _T_332;
  wire  _T_334;
  wire  _T_336;
  wire  _T_338;
  wire  _T_340;
  wire  _T_342;
  wire  _T_344;
  wire  _T_347_0;
  wire  _T_347_1;
  wire  _T_347_2;
  wire  _T_347_3;
  wire  _T_347_4;
  wire  _T_357;
  wire  _T_359;
  wire  _T_361;
  wire  _T_363;
  wire  _T_365;
  wire  _T_366;
  wire  _T_367;
  wire  _T_368;
  wire  _T_369;
  wire  _T_371;
  wire  _T_373;
  wire  _T_375;
  wire  _T_377;
  wire  _T_379;
  wire  _T_381;
  wire  _T_384_0;
  wire  _T_384_1;
  wire  _T_384_2;
  wire  _T_384_3;
  wire  _T_384_4;
  wire  _T_394;
  wire  _T_396;
  wire  _T_398;
  wire  _T_400;
  wire  _T_402;
  wire  _T_403;
  wire  _T_404;
  wire  _T_405;
  wire  _T_406;
  wire  _T_408;
  FF_103 ff_0 (
    .clock(ff_0_clock),
    .reset(ff_0_reset),
    .io_input_0_data(ff_0_io_input_0_data),
    .io_input_0_enable(ff_0_io_input_0_enable),
    .io_input_0_reset(ff_0_io_input_0_reset),
    .io_output_data(ff_0_io_output_data)
  );
  FF_103 ff_1 (
    .clock(ff_1_clock),
    .reset(ff_1_reset),
    .io_input_0_data(ff_1_io_input_0_data),
    .io_input_0_enable(ff_1_io_input_0_enable),
    .io_input_0_reset(ff_1_io_input_0_reset),
    .io_output_data(ff_1_io_output_data)
  );
  FF_103 ff_2 (
    .clock(ff_2_clock),
    .reset(ff_2_reset),
    .io_input_0_data(ff_2_io_input_0_data),
    .io_input_0_enable(ff_2_io_input_0_enable),
    .io_input_0_reset(ff_2_io_input_0_reset),
    .io_output_data(ff_2_io_output_data)
  );
  FF_103 ff_3 (
    .clock(ff_3_clock),
    .reset(ff_3_reset),
    .io_input_0_data(ff_3_io_input_0_data),
    .io_input_0_enable(ff_3_io_input_0_enable),
    .io_input_0_reset(ff_3_io_input_0_reset),
    .io_output_data(ff_3_io_output_data)
  );
  FF_103 ff_4 (
    .clock(ff_4_clock),
    .reset(ff_4_reset),
    .io_input_0_data(ff_4_io_input_0_data),
    .io_input_0_enable(ff_4_io_input_0_enable),
    .io_input_0_reset(ff_4_io_input_0_reset),
    .io_output_data(ff_4_io_output_data)
  );
  SRFF sEn_latch_0 (
    .clock(sEn_latch_0_clock),
    .reset(sEn_latch_0_reset),
    .io_input_set(sEn_latch_0_io_input_set),
    .io_input_reset(sEn_latch_0_io_input_reset),
    .io_input_asyn_reset(sEn_latch_0_io_input_asyn_reset),
    .io_output_data(sEn_latch_0_io_output_data)
  );
  SRFF sEn_latch_1 (
    .clock(sEn_latch_1_clock),
    .reset(sEn_latch_1_reset),
    .io_input_set(sEn_latch_1_io_input_set),
    .io_input_reset(sEn_latch_1_io_input_reset),
    .io_input_asyn_reset(sEn_latch_1_io_input_asyn_reset),
    .io_output_data(sEn_latch_1_io_output_data)
  );
  SRFF sEn_latch_2 (
    .clock(sEn_latch_2_clock),
    .reset(sEn_latch_2_reset),
    .io_input_set(sEn_latch_2_io_input_set),
    .io_input_reset(sEn_latch_2_io_input_reset),
    .io_input_asyn_reset(sEn_latch_2_io_input_asyn_reset),
    .io_output_data(sEn_latch_2_io_output_data)
  );
  SRFF sEn_latch_3 (
    .clock(sEn_latch_3_clock),
    .reset(sEn_latch_3_reset),
    .io_input_set(sEn_latch_3_io_input_set),
    .io_input_reset(sEn_latch_3_io_input_reset),
    .io_input_asyn_reset(sEn_latch_3_io_input_asyn_reset),
    .io_output_data(sEn_latch_3_io_output_data)
  );
  SRFF sEn_latch_4 (
    .clock(sEn_latch_4_clock),
    .reset(sEn_latch_4_reset),
    .io_input_set(sEn_latch_4_io_input_set),
    .io_input_reset(sEn_latch_4_io_input_reset),
    .io_input_asyn_reset(sEn_latch_4_io_input_asyn_reset),
    .io_output_data(sEn_latch_4_io_output_data)
  );
  SRFF sDone_latch_0 (
    .clock(sDone_latch_0_clock),
    .reset(sDone_latch_0_reset),
    .io_input_set(sDone_latch_0_io_input_set),
    .io_input_reset(sDone_latch_0_io_input_reset),
    .io_input_asyn_reset(sDone_latch_0_io_input_asyn_reset),
    .io_output_data(sDone_latch_0_io_output_data)
  );
  SRFF sDone_latch_1 (
    .clock(sDone_latch_1_clock),
    .reset(sDone_latch_1_reset),
    .io_input_set(sDone_latch_1_io_input_set),
    .io_input_reset(sDone_latch_1_io_input_reset),
    .io_input_asyn_reset(sDone_latch_1_io_input_asyn_reset),
    .io_output_data(sDone_latch_1_io_output_data)
  );
  SRFF sDone_latch_2 (
    .clock(sDone_latch_2_clock),
    .reset(sDone_latch_2_reset),
    .io_input_set(sDone_latch_2_io_input_set),
    .io_input_reset(sDone_latch_2_io_input_reset),
    .io_input_asyn_reset(sDone_latch_2_io_input_asyn_reset),
    .io_output_data(sDone_latch_2_io_output_data)
  );
  SRFF sDone_latch_3 (
    .clock(sDone_latch_3_clock),
    .reset(sDone_latch_3_reset),
    .io_input_set(sDone_latch_3_io_input_set),
    .io_input_reset(sDone_latch_3_io_input_reset),
    .io_input_asyn_reset(sDone_latch_3_io_input_asyn_reset),
    .io_output_data(sDone_latch_3_io_output_data)
  );
  SRFF sDone_latch_4 (
    .clock(sDone_latch_4_clock),
    .reset(sDone_latch_4_reset),
    .io_input_set(sDone_latch_4_io_input_set),
    .io_input_reset(sDone_latch_4_io_input_reset),
    .io_input_asyn_reset(sDone_latch_4_io_input_asyn_reset),
    .io_output_data(sDone_latch_4_io_output_data)
  );
  RetimeWrapper RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 (
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 (
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 (
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 (
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 (
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 (
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 (
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper RetimeWrapper_8 (
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper RetimeWrapper_9 (
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper RetimeWrapper_10 (
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper RetimeWrapper_11 (
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper RetimeWrapper_12 (
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper RetimeWrapper_13 (
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper RetimeWrapper_14 (
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper RetimeWrapper_15 (
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper RetimeWrapper_16 (
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper RetimeWrapper_17 (
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper RetimeWrapper_18 (
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper RetimeWrapper_19 (
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper RetimeWrapper_20 (
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper RetimeWrapper_21 (
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper RetimeWrapper_22 (
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper RetimeWrapper_23 (
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper RetimeWrapper_24 (
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  NBufCtr statesIn_0 (
    .clock(statesIn_0_clock),
    .reset(statesIn_0_reset),
    .io_input_enable(statesIn_0_io_input_enable),
    .io_output_count(statesIn_0_io_output_count)
  );
  NBufCtr_1 statesOut_0 (
    .clock(statesOut_0_clock),
    .reset(statesOut_0_reset),
    .io_input_enable(statesOut_0_io_input_enable)
  );
  NBufCtr_2 statesOut_1 (
    .clock(statesOut_1_clock),
    .reset(statesOut_1_reset),
    .io_input_enable(statesOut_1_io_input_enable),
    .io_output_count(statesOut_1_io_output_count)
  );
  NBufCtr_3 statesOut_2 (
    .clock(statesOut_2_clock),
    .reset(statesOut_2_reset),
    .io_input_enable(statesOut_2_io_input_enable),
    .io_output_count(statesOut_2_io_output_count)
  );
  NBufCtr_4 statesOut_3 (
    .clock(statesOut_3_clock),
    .reset(statesOut_3_reset),
    .io_input_enable(statesOut_3_io_input_enable),
    .io_output_count(statesOut_3_io_output_count)
  );
  NBufCtr_5 statesOut_4 (
    .clock(statesOut_4_clock),
    .reset(statesOut_4_reset),
    .io_input_enable(statesOut_4_io_input_enable),
    .io_output_count(statesOut_4_io_output_count)
  );
  assign _T_20 = ~ io_sDone_0;
  assign _T_21 = io_sEn_0 & _T_20;
  assign _T_22 = io_sEn_0 & io_sDone_0;
  assign _T_23 = ~ io_sEn_0;
  assign _T_28 = _T_22 & _T_27;
  assign _T_29 = _T_21 | _T_28;
  assign _T_34 = swap | _T_33;
  assign _T_43 = swap | _T_42;
  assign _T_48 = ~ io_sDone_1;
  assign _T_49 = io_sEn_1 & _T_48;
  assign _T_50 = io_sEn_1 & io_sDone_1;
  assign _T_51 = ~ io_sEn_1;
  assign _T_56 = _T_50 & _T_55;
  assign _T_57 = _T_49 | _T_56;
  assign _T_62 = swap | _T_61;
  assign _T_71 = swap | _T_70;
  assign _T_76 = ~ io_sDone_2;
  assign _T_77 = io_sEn_2 & _T_76;
  assign _T_78 = io_sEn_2 & io_sDone_2;
  assign _T_79 = ~ io_sEn_2;
  assign _T_84 = _T_78 & _T_83;
  assign _T_85 = _T_77 | _T_84;
  assign _T_90 = swap | _T_89;
  assign _T_99 = swap | _T_98;
  assign _T_104 = ~ io_sDone_3;
  assign _T_105 = io_sEn_3 & _T_104;
  assign _T_106 = io_sEn_3 & io_sDone_3;
  assign _T_107 = ~ io_sEn_3;
  assign _T_112 = _T_106 & _T_111;
  assign _T_113 = _T_105 | _T_112;
  assign _T_118 = swap | _T_117;
  assign _T_127 = swap | _T_126;
  assign _T_132 = ~ io_sDone_4;
  assign _T_133 = io_sEn_4 & _T_132;
  assign _T_134 = io_sEn_4 & io_sDone_4;
  assign _T_135 = ~ io_sEn_4;
  assign _T_140 = _T_134 & _T_139;
  assign _T_141 = _T_133 | _T_140;
  assign _T_146 = swap | _T_145;
  assign _T_155 = swap | _T_154;
  assign _T_160 = sEn_latch_0_io_output_data | sEn_latch_1_io_output_data;
  assign _T_161 = _T_160 | sEn_latch_2_io_output_data;
  assign _T_162 = _T_161 | sEn_latch_3_io_output_data;
  assign anyEnabled = _T_162 | sEn_latch_4_io_output_data;
  assign _T_163 = sDone_latch_0_io_output_data | io_sDone_0;
  assign _T_164 = sEn_latch_0_io_output_data == _T_163;
  assign _T_165 = sDone_latch_1_io_output_data | io_sDone_1;
  assign _T_166 = sEn_latch_1_io_output_data == _T_165;
  assign _T_167 = sDone_latch_2_io_output_data | io_sDone_2;
  assign _T_168 = sEn_latch_2_io_output_data == _T_167;
  assign _T_169 = sDone_latch_3_io_output_data | io_sDone_3;
  assign _T_170 = sEn_latch_3_io_output_data == _T_169;
  assign _T_171 = sDone_latch_4_io_output_data | io_sDone_4;
  assign _T_172 = sEn_latch_4_io_output_data == _T_171;
  assign _T_173 = _T_164 & _T_166;
  assign _T_174 = _T_173 & _T_168;
  assign _T_175 = _T_174 & _T_170;
  assign _T_176 = _T_175 & _T_172;
  assign _T_177 = _T_176 & anyEnabled;
  assign _T_178 = ~ _T_177;
  assign _T_187 = _T_177 & _T_181;
  assign _T_195 = statesIn_0_io_output_count == 4'h0;
  assign _T_198 = io_input_0_enable & _T_195;
  assign _T_201 = statesIn_0_io_output_count == 4'h1;
  assign _T_204 = io_input_0_enable & _T_201;
  assign _T_207 = statesIn_0_io_output_count == 4'h2;
  assign _T_210 = io_input_0_enable & _T_207;
  assign _T_213 = statesIn_0_io_output_count == 4'h3;
  assign _T_216 = io_input_0_enable & _T_213;
  assign _T_219 = statesIn_0_io_output_count == 4'h4;
  assign _T_222 = io_input_0_enable & _T_219;
  assign _T_262 = statesOut_1_io_output_count == 4'h0;
  assign _T_264 = statesOut_1_io_output_count == 4'h1;
  assign _T_266 = statesOut_1_io_output_count == 4'h2;
  assign _T_268 = statesOut_1_io_output_count == 4'h3;
  assign _T_270 = statesOut_1_io_output_count == 4'h4;
  assign _T_283 = _T_262 ? _T_273_0 : 1'h0;
  assign _T_285 = _T_264 ? _T_273_1 : 1'h0;
  assign _T_287 = _T_266 ? _T_273_2 : 1'h0;
  assign _T_289 = _T_268 ? _T_273_3 : 1'h0;
  assign _T_291 = _T_270 ? _T_273_4 : 1'h0;
  assign _T_292 = _T_283 | _T_285;
  assign _T_293 = _T_292 | _T_287;
  assign _T_294 = _T_293 | _T_289;
  assign _T_295 = _T_294 | _T_291;
  assign _T_299 = statesOut_2_io_output_count == 4'h0;
  assign _T_301 = statesOut_2_io_output_count == 4'h1;
  assign _T_303 = statesOut_2_io_output_count == 4'h2;
  assign _T_305 = statesOut_2_io_output_count == 4'h3;
  assign _T_307 = statesOut_2_io_output_count == 4'h4;
  assign _T_320 = _T_299 ? _T_310_0 : 1'h0;
  assign _T_322 = _T_301 ? _T_310_1 : 1'h0;
  assign _T_324 = _T_303 ? _T_310_2 : 1'h0;
  assign _T_326 = _T_305 ? _T_310_3 : 1'h0;
  assign _T_328 = _T_307 ? _T_310_4 : 1'h0;
  assign _T_329 = _T_320 | _T_322;
  assign _T_330 = _T_329 | _T_324;
  assign _T_331 = _T_330 | _T_326;
  assign _T_332 = _T_331 | _T_328;
  assign _T_336 = statesOut_3_io_output_count == 4'h0;
  assign _T_338 = statesOut_3_io_output_count == 4'h1;
  assign _T_340 = statesOut_3_io_output_count == 4'h2;
  assign _T_342 = statesOut_3_io_output_count == 4'h3;
  assign _T_344 = statesOut_3_io_output_count == 4'h4;
  assign _T_357 = _T_336 ? _T_347_0 : 1'h0;
  assign _T_359 = _T_338 ? _T_347_1 : 1'h0;
  assign _T_361 = _T_340 ? _T_347_2 : 1'h0;
  assign _T_363 = _T_342 ? _T_347_3 : 1'h0;
  assign _T_365 = _T_344 ? _T_347_4 : 1'h0;
  assign _T_366 = _T_357 | _T_359;
  assign _T_367 = _T_366 | _T_361;
  assign _T_368 = _T_367 | _T_363;
  assign _T_369 = _T_368 | _T_365;
  assign _T_373 = statesOut_4_io_output_count == 4'h0;
  assign _T_375 = statesOut_4_io_output_count == 4'h1;
  assign _T_377 = statesOut_4_io_output_count == 4'h2;
  assign _T_379 = statesOut_4_io_output_count == 4'h3;
  assign _T_381 = statesOut_4_io_output_count == 4'h4;
  assign _T_394 = _T_373 ? _T_384_0 : 1'h0;
  assign _T_396 = _T_375 ? _T_384_1 : 1'h0;
  assign _T_398 = _T_377 ? _T_384_2 : 1'h0;
  assign _T_400 = _T_379 ? _T_384_3 : 1'h0;
  assign _T_402 = _T_381 ? _T_384_4 : 1'h0;
  assign _T_403 = _T_394 | _T_396;
  assign _T_404 = _T_403 | _T_398;
  assign _T_405 = _T_404 | _T_400;
  assign _T_406 = _T_405 | _T_402;
  assign io_output_1_data = _T_297;
  assign io_output_2_data = _T_334;
  assign io_output_3_data = _T_371;
  assign io_output_4_data = _T_408;
  assign ff_0_io_input_0_data = _T_197_data;
  assign ff_0_io_input_0_enable = _T_197_enable;
  assign ff_0_io_input_0_reset = _T_197_reset;
  assign ff_0_clock = clock;
  assign ff_0_reset = reset;
  assign ff_1_io_input_0_data = _T_203_data;
  assign ff_1_io_input_0_enable = _T_203_enable;
  assign ff_1_io_input_0_reset = _T_203_reset;
  assign ff_1_clock = clock;
  assign ff_1_reset = reset;
  assign ff_2_io_input_0_data = _T_209_data;
  assign ff_2_io_input_0_enable = _T_209_enable;
  assign ff_2_io_input_0_reset = _T_209_reset;
  assign ff_2_clock = clock;
  assign ff_2_reset = reset;
  assign ff_3_io_input_0_data = _T_215_data;
  assign ff_3_io_input_0_enable = _T_215_enable;
  assign ff_3_io_input_0_reset = _T_215_reset;
  assign ff_3_clock = clock;
  assign ff_3_reset = reset;
  assign ff_4_io_input_0_data = _T_221_data;
  assign ff_4_io_input_0_enable = _T_221_enable;
  assign ff_4_io_input_0_reset = _T_221_reset;
  assign ff_4_clock = clock;
  assign ff_4_reset = reset;
  assign sEn_latch_0_io_input_set = _T_29;
  assign sEn_latch_0_io_input_reset = _T_34;
  assign sEn_latch_0_io_input_asyn_reset = _T_38;
  assign sEn_latch_0_clock = clock;
  assign sEn_latch_0_reset = reset;
  assign sEn_latch_1_io_input_set = _T_57;
  assign sEn_latch_1_io_input_reset = _T_62;
  assign sEn_latch_1_io_input_asyn_reset = _T_66;
  assign sEn_latch_1_clock = clock;
  assign sEn_latch_1_reset = reset;
  assign sEn_latch_2_io_input_set = _T_85;
  assign sEn_latch_2_io_input_reset = _T_90;
  assign sEn_latch_2_io_input_asyn_reset = _T_94;
  assign sEn_latch_2_clock = clock;
  assign sEn_latch_2_reset = reset;
  assign sEn_latch_3_io_input_set = _T_113;
  assign sEn_latch_3_io_input_reset = _T_118;
  assign sEn_latch_3_io_input_asyn_reset = _T_122;
  assign sEn_latch_3_clock = clock;
  assign sEn_latch_3_reset = reset;
  assign sEn_latch_4_io_input_set = _T_141;
  assign sEn_latch_4_io_input_reset = _T_146;
  assign sEn_latch_4_io_input_asyn_reset = _T_150;
  assign sEn_latch_4_clock = clock;
  assign sEn_latch_4_reset = reset;
  assign sDone_latch_0_io_input_set = io_sDone_0;
  assign sDone_latch_0_io_input_reset = _T_43;
  assign sDone_latch_0_io_input_asyn_reset = _T_47;
  assign sDone_latch_0_clock = clock;
  assign sDone_latch_0_reset = reset;
  assign sDone_latch_1_io_input_set = io_sDone_1;
  assign sDone_latch_1_io_input_reset = _T_71;
  assign sDone_latch_1_io_input_asyn_reset = _T_75;
  assign sDone_latch_1_clock = clock;
  assign sDone_latch_1_reset = reset;
  assign sDone_latch_2_io_input_set = io_sDone_2;
  assign sDone_latch_2_io_input_reset = _T_99;
  assign sDone_latch_2_io_input_asyn_reset = _T_103;
  assign sDone_latch_2_clock = clock;
  assign sDone_latch_2_reset = reset;
  assign sDone_latch_3_io_input_set = io_sDone_3;
  assign sDone_latch_3_io_input_reset = _T_127;
  assign sDone_latch_3_io_input_asyn_reset = _T_131;
  assign sDone_latch_3_clock = clock;
  assign sDone_latch_3_reset = reset;
  assign sDone_latch_4_io_input_set = io_sDone_4;
  assign sDone_latch_4_io_input_reset = _T_155;
  assign sDone_latch_4_io_input_asyn_reset = _T_159;
  assign sDone_latch_4_clock = clock;
  assign sDone_latch_4_reset = reset;
  assign swap = _T_187;
  assign RetimeWrapper_io_flow = 1'h1;
  assign RetimeWrapper_io_in = _T_23;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_27 = RetimeWrapper_io_out;
  assign RetimeWrapper_1_io_flow = 1'h1;
  assign RetimeWrapper_1_io_in = swap;
  assign RetimeWrapper_1_clock = clock;
  assign RetimeWrapper_1_reset = reset;
  assign _T_33 = RetimeWrapper_1_io_out;
  assign RetimeWrapper_2_io_flow = 1'h1;
  assign RetimeWrapper_2_io_in = reset;
  assign RetimeWrapper_2_clock = clock;
  assign RetimeWrapper_2_reset = reset;
  assign _T_38 = RetimeWrapper_2_io_out;
  assign RetimeWrapper_3_io_flow = 1'h1;
  assign RetimeWrapper_3_io_in = swap;
  assign RetimeWrapper_3_clock = clock;
  assign RetimeWrapper_3_reset = reset;
  assign _T_42 = RetimeWrapper_3_io_out;
  assign RetimeWrapper_4_io_flow = 1'h1;
  assign RetimeWrapper_4_io_in = reset;
  assign RetimeWrapper_4_clock = clock;
  assign RetimeWrapper_4_reset = reset;
  assign _T_47 = RetimeWrapper_4_io_out;
  assign RetimeWrapper_5_io_flow = 1'h1;
  assign RetimeWrapper_5_io_in = _T_51;
  assign RetimeWrapper_5_clock = clock;
  assign RetimeWrapper_5_reset = reset;
  assign _T_55 = RetimeWrapper_5_io_out;
  assign RetimeWrapper_6_io_flow = 1'h1;
  assign RetimeWrapper_6_io_in = swap;
  assign RetimeWrapper_6_clock = clock;
  assign RetimeWrapper_6_reset = reset;
  assign _T_61 = RetimeWrapper_6_io_out;
  assign RetimeWrapper_7_io_flow = 1'h1;
  assign RetimeWrapper_7_io_in = reset;
  assign RetimeWrapper_7_clock = clock;
  assign RetimeWrapper_7_reset = reset;
  assign _T_66 = RetimeWrapper_7_io_out;
  assign RetimeWrapper_8_io_flow = 1'h1;
  assign RetimeWrapper_8_io_in = swap;
  assign RetimeWrapper_8_clock = clock;
  assign RetimeWrapper_8_reset = reset;
  assign _T_70 = RetimeWrapper_8_io_out;
  assign RetimeWrapper_9_io_flow = 1'h1;
  assign RetimeWrapper_9_io_in = reset;
  assign RetimeWrapper_9_clock = clock;
  assign RetimeWrapper_9_reset = reset;
  assign _T_75 = RetimeWrapper_9_io_out;
  assign RetimeWrapper_10_io_flow = 1'h1;
  assign RetimeWrapper_10_io_in = _T_79;
  assign RetimeWrapper_10_clock = clock;
  assign RetimeWrapper_10_reset = reset;
  assign _T_83 = RetimeWrapper_10_io_out;
  assign RetimeWrapper_11_io_flow = 1'h1;
  assign RetimeWrapper_11_io_in = swap;
  assign RetimeWrapper_11_clock = clock;
  assign RetimeWrapper_11_reset = reset;
  assign _T_89 = RetimeWrapper_11_io_out;
  assign RetimeWrapper_12_io_flow = 1'h1;
  assign RetimeWrapper_12_io_in = reset;
  assign RetimeWrapper_12_clock = clock;
  assign RetimeWrapper_12_reset = reset;
  assign _T_94 = RetimeWrapper_12_io_out;
  assign RetimeWrapper_13_io_flow = 1'h1;
  assign RetimeWrapper_13_io_in = swap;
  assign RetimeWrapper_13_clock = clock;
  assign RetimeWrapper_13_reset = reset;
  assign _T_98 = RetimeWrapper_13_io_out;
  assign RetimeWrapper_14_io_flow = 1'h1;
  assign RetimeWrapper_14_io_in = reset;
  assign RetimeWrapper_14_clock = clock;
  assign RetimeWrapper_14_reset = reset;
  assign _T_103 = RetimeWrapper_14_io_out;
  assign RetimeWrapper_15_io_flow = 1'h1;
  assign RetimeWrapper_15_io_in = _T_107;
  assign RetimeWrapper_15_clock = clock;
  assign RetimeWrapper_15_reset = reset;
  assign _T_111 = RetimeWrapper_15_io_out;
  assign RetimeWrapper_16_io_flow = 1'h1;
  assign RetimeWrapper_16_io_in = swap;
  assign RetimeWrapper_16_clock = clock;
  assign RetimeWrapper_16_reset = reset;
  assign _T_117 = RetimeWrapper_16_io_out;
  assign RetimeWrapper_17_io_flow = 1'h1;
  assign RetimeWrapper_17_io_in = reset;
  assign RetimeWrapper_17_clock = clock;
  assign RetimeWrapper_17_reset = reset;
  assign _T_122 = RetimeWrapper_17_io_out;
  assign RetimeWrapper_18_io_flow = 1'h1;
  assign RetimeWrapper_18_io_in = swap;
  assign RetimeWrapper_18_clock = clock;
  assign RetimeWrapper_18_reset = reset;
  assign _T_126 = RetimeWrapper_18_io_out;
  assign RetimeWrapper_19_io_flow = 1'h1;
  assign RetimeWrapper_19_io_in = reset;
  assign RetimeWrapper_19_clock = clock;
  assign RetimeWrapper_19_reset = reset;
  assign _T_131 = RetimeWrapper_19_io_out;
  assign RetimeWrapper_20_io_flow = 1'h1;
  assign RetimeWrapper_20_io_in = _T_135;
  assign RetimeWrapper_20_clock = clock;
  assign RetimeWrapper_20_reset = reset;
  assign _T_139 = RetimeWrapper_20_io_out;
  assign RetimeWrapper_21_io_flow = 1'h1;
  assign RetimeWrapper_21_io_in = swap;
  assign RetimeWrapper_21_clock = clock;
  assign RetimeWrapper_21_reset = reset;
  assign _T_145 = RetimeWrapper_21_io_out;
  assign RetimeWrapper_22_io_flow = 1'h1;
  assign RetimeWrapper_22_io_in = reset;
  assign RetimeWrapper_22_clock = clock;
  assign RetimeWrapper_22_reset = reset;
  assign _T_150 = RetimeWrapper_22_io_out;
  assign RetimeWrapper_23_io_flow = 1'h1;
  assign RetimeWrapper_23_io_in = swap;
  assign RetimeWrapper_23_clock = clock;
  assign RetimeWrapper_23_reset = reset;
  assign _T_154 = RetimeWrapper_23_io_out;
  assign RetimeWrapper_24_io_flow = 1'h1;
  assign RetimeWrapper_24_io_in = reset;
  assign RetimeWrapper_24_clock = clock;
  assign RetimeWrapper_24_reset = reset;
  assign _T_159 = RetimeWrapper_24_io_out;
  assign statesIn_0_io_input_enable = swap;
  assign statesIn_0_clock = clock;
  assign statesIn_0_reset = reset;
  assign statesOut_0_io_input_enable = swap;
  assign statesOut_0_clock = clock;
  assign statesOut_0_reset = reset;
  assign statesOut_1_io_input_enable = swap;
  assign statesOut_1_clock = clock;
  assign statesOut_1_reset = reset;
  assign statesOut_2_io_input_enable = swap;
  assign statesOut_2_clock = clock;
  assign statesOut_2_reset = reset;
  assign statesOut_3_io_input_enable = swap;
  assign statesOut_3_clock = clock;
  assign statesOut_3_reset = reset;
  assign statesOut_4_io_input_enable = swap;
  assign statesOut_4_clock = clock;
  assign statesOut_4_reset = reset;
  assign _T_197_data = io_input_0_data;
  assign _T_197_enable = _T_198;
  assign _T_197_reset = io_input_0_reset;
  assign _T_203_data = io_input_0_data;
  assign _T_203_enable = _T_204;
  assign _T_203_reset = io_input_0_reset;
  assign _T_209_data = io_input_0_data;
  assign _T_209_enable = _T_210;
  assign _T_209_reset = io_input_0_reset;
  assign _T_215_data = io_input_0_data;
  assign _T_215_enable = _T_216;
  assign _T_215_reset = io_input_0_reset;
  assign _T_221_data = io_input_0_data;
  assign _T_221_enable = _T_222;
  assign _T_221_reset = io_input_0_reset;
  assign _T_273_0 = ff_0_io_output_data;
  assign _T_273_1 = ff_1_io_output_data;
  assign _T_273_2 = ff_2_io_output_data;
  assign _T_273_3 = ff_3_io_output_data;
  assign _T_273_4 = ff_4_io_output_data;
  assign _T_297 = _T_295;
  assign _T_310_0 = ff_0_io_output_data;
  assign _T_310_1 = ff_1_io_output_data;
  assign _T_310_2 = ff_2_io_output_data;
  assign _T_310_3 = ff_3_io_output_data;
  assign _T_310_4 = ff_4_io_output_data;
  assign _T_334 = _T_332;
  assign _T_347_0 = ff_0_io_output_data;
  assign _T_347_1 = ff_1_io_output_data;
  assign _T_347_2 = ff_2_io_output_data;
  assign _T_347_3 = ff_3_io_output_data;
  assign _T_347_4 = ff_4_io_output_data;
  assign _T_371 = _T_369;
  assign _T_384_0 = ff_0_io_output_data;
  assign _T_384_1 = ff_1_io_output_data;
  assign _T_384_2 = ff_2_io_output_data;
  assign _T_384_3 = ff_3_io_output_data;
  assign _T_384_4 = ff_4_io_output_data;
  assign _T_408 = _T_406;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_181 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_181 <= 1'h0;
    end else begin
      _T_181 <= _T_178;
    end
  end
endmodule
module SingleCounter_19(
  input   clock,
  input   reset,
  input   io_input_reset,
  output  io_output_done
);
  wire  FF_clock;
  wire  FF_reset;
  wire [31:0] FF_io_input_0_data;
  wire [31:0] FF_io_input_0_init;
  wire  FF_io_input_0_enable;
  wire  FF_io_input_0_reset;
  wire [31:0] FF_io_output_data;
  wire [31:0] _T_21;
  wire [32:0] _T_23;
  wire [31:0] _T_24;
  wire [31:0] _T_25;
  wire  _T_29;
  wire [31:0] _T_40;
  wire [31:0] _T_43;
  wire [31:0] _T_44;
  wire [31:0] _T_45;
  FF_1 FF (
    .clock(FF_clock),
    .reset(FF_reset),
    .io_input_0_data(FF_io_input_0_data),
    .io_input_0_init(FF_io_input_0_init),
    .io_input_0_enable(FF_io_input_0_enable),
    .io_input_0_reset(FF_io_input_0_reset),
    .io_output_data(FF_io_output_data)
  );
  assign _T_21 = $signed(FF_io_output_data);
  assign _T_23 = $signed(_T_21) + $signed(32'sh1);
  assign _T_24 = _T_23[31:0];
  assign _T_25 = $signed(_T_24);
  assign _T_29 = $signed(_T_25) >= $signed(32'sh6);
  assign _T_40 = $unsigned(_T_21);
  assign _T_43 = $unsigned(_T_25);
  assign _T_44 = _T_29 ? _T_40 : _T_43;
  assign _T_45 = io_input_reset ? 32'h0 : _T_44;
  assign io_output_done = _T_29;
  assign FF_io_input_0_data = _T_45;
  assign FF_io_input_0_init = 32'h0;
  assign FF_io_input_0_enable = 1'h1;
  assign FF_io_input_0_reset = io_input_reset;
  assign FF_clock = clock;
  assign FF_reset = reset;
endmodule
module AccelTop(
  input         clock,
  input         reset,
  input         io_enable,
  output        io_done,
  input         io_memStreams_loads_3_cmd_ready,
  output        io_memStreams_loads_3_cmd_valid,
  output [63:0] io_memStreams_loads_3_cmd_bits_addr,
  output        io_memStreams_loads_3_cmd_bits_isWr,
  output [15:0] io_memStreams_loads_3_cmd_bits_size,
  output        io_memStreams_loads_3_rdata_ready,
  input         io_memStreams_loads_3_rdata_valid,
  input  [31:0] io_memStreams_loads_3_rdata_bits_0,
  input         io_memStreams_loads_2_cmd_ready,
  output        io_memStreams_loads_2_cmd_valid,
  output [63:0] io_memStreams_loads_2_cmd_bits_addr,
  output        io_memStreams_loads_2_cmd_bits_isWr,
  output [15:0] io_memStreams_loads_2_cmd_bits_size,
  output        io_memStreams_loads_2_rdata_ready,
  input         io_memStreams_loads_2_rdata_valid,
  input  [31:0] io_memStreams_loads_2_rdata_bits_0,
  input         io_memStreams_loads_1_cmd_ready,
  output        io_memStreams_loads_1_cmd_valid,
  output [63:0] io_memStreams_loads_1_cmd_bits_addr,
  output        io_memStreams_loads_1_cmd_bits_isWr,
  output [15:0] io_memStreams_loads_1_cmd_bits_size,
  output        io_memStreams_loads_1_rdata_ready,
  input         io_memStreams_loads_1_rdata_valid,
  input  [31:0] io_memStreams_loads_1_rdata_bits_0,
  input         io_memStreams_loads_0_cmd_ready,
  output        io_memStreams_loads_0_cmd_valid,
  output [63:0] io_memStreams_loads_0_cmd_bits_addr,
  output        io_memStreams_loads_0_cmd_bits_isWr,
  output [15:0] io_memStreams_loads_0_cmd_bits_size,
  output        io_memStreams_loads_0_rdata_ready,
  input         io_memStreams_loads_0_rdata_valid,
  input  [31:0] io_memStreams_loads_0_rdata_bits_0,
  input  [63:0] io_argIns_0,
  input  [63:0] io_argIns_1,
  input  [63:0] io_argIns_2,
  output        io_argOuts_0_valid,
  output [63:0] io_argOuts_0_bits
);
  wire [63:0] x3141_data_options_0;
  wire  x3141_en_options_0;
  wire  RootController_done;
  wire  RootController_en;
  wire  RootController_resetter;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire  RetimeWrapper_io_flow;
  wire  RetimeWrapper_io_in;
  wire  RetimeWrapper_io_out;
  wire  retime_released;
  wire [31:0] x3153_number;
  wire  x3155_en;
  wire  x3155_resetter;
  wire [31:0] x3154_0;
  wire [31:0] x3154_1;
  wire [31:0] x3515_level0_iters;
  wire  x3515_done;
  wire  x3515_en;
  wire  x3515_base_en;
  wire  x3515_resetter;
  wire  x3515_ctr_trivial;
  wire  x3515_rst_en;
  wire  x3152_wren;
  wire  x3152_resetter;
  wire [31:0] b1202_number;
  wire [31:0] b1203_number;
  wire  x3174_done;
  wire  x3174_en;
  wire  x3174_base_en;
  wire  x3174_resetter;
  wire  x3174_ctr_trivial;
  wire  x3167_done;
  wire  x3167_en;
  wire  x3167_base_en;
  wire  x3167_mask;
  wire  x3167_resetter;
  wire  x3167_datapath_en;
  wire  x3167_ctr_trivial;
  wire [31:0] x3162_number;
  wire [31:0] x3163_number;
  wire [31:0] x3164_number;
  wire  x3173_done;
  wire  x3173_en;
  wire  x3173_base_en;
  wire  x3173_mask;
  wire  x3173_resetter;
  wire  x3173_datapath_en;
  wire  x3173_ctr_trivial;
  wire [31:0] x3168_number;
  wire [31:0] x3169_number;
  wire [31:0] x3170_number;
  wire  x3301_done;
  wire  x3301_en;
  wire  x3301_base_en;
  wire  x3301_resetter;
  wire  x3301_ctr_trivial;
  wire  x3237_done;
  wire  x3237_en;
  wire  x3237_base_en;
  wire  x3237_mask;
  wire  x3237_resetter;
  wire  x3237_ctr_trivial;
  wire  x3175_valid_options_0;
  wire  x3175_valid_stops_0;
  wire  x3175_valid;
  wire [96:0] x3175_data_options_0;
  wire  x3175_ready;
  wire  x3177_ready_options_0;
  wire  x3177_ready;
  wire  x3177_now_valid;
  wire  x3177_valid;
  wire [31:0] x3177_0_number;
  wire  x3208_done;
  wire  x3208_en;
  wire  x3208_base_en;
  wire  x3208_mask;
  wire  x3208_resetter;
  wire  x3208_datapath_en;
  wire  x3208_ctr_trivial;
  wire [31:0] x3178_number;
  wire [31:0] x3179_number;
  wire [31:0] x3182_number;
  wire [31:0] x3183_number;
  wire [31:0] x3184_number;
  wire [31:0] x3185_number;
  wire [31:0] x3186_number;
  wire [31:0] x3189_number;
  wire  x3190;
  wire [31:0] x3191_number;
  wire [31:0] x3192_number;
  wire [31:0] x3193_number;
  wire [31:0] x3194_number;
  wire [31:0] x3195_number;
  wire [31:0] x3196_number;
  wire [31:0] x3197_number;
  wire [31:0] x3198_number;
  wire [31:0] x3199_number;
  wire [63:0] x3200_number;
  wire [63:0] x3202_number;
  wire [63:0] x3203_number;
  wire [63:0] x3204_item0;
  wire [31:0] x3204_item1;
  wire [96:0] x3204;
  wire [31:0] x3206_item0;
  wire [31:0] x3206_item1;
  wire [31:0] x3206_item2;
  wire [95:0] x3206;
  wire  x3236_done;
  wire  x3236_en;
  wire  x3236_base_en;
  wire  x3236_mask;
  wire  x3236_resetter;
  wire  x3236_ctr_trivial;
  wire  x3220_done;
  wire  x3220_en;
  wire  x3220_base_en;
  wire  x3220_mask;
  wire  x3220_resetter;
  wire  x3220_datapath_en;
  wire  x3220_ctr_trivial;
  wire [31:0] x3214_number;
  wire [31:0] x3216_number;
  wire [31:0] x3218_number;
  wire [31:0] x3221_number;
  wire  x3223_done;
  wire  x3223_en;
  wire  x3223_resetter;
  wire [31:0] x3222_0;
  wire  x3235_done;
  wire  x3235_en;
  wire  x3235_base_en;
  wire  x3235_mask;
  wire  x3235_datapath_en;
  wire  x3235_ctr_trivial;
  wire [31:0] b1270_number;
  wire [31:0] x3224_number;
  wire  x3225;
  wire [31:0] x3226_number;
  wire  x3227;
  wire  x3228;
  wire [31:0] x3229_number;
  wire  x3230;
  wire [31:0] x3232_number;
  wire  x3233;
  wire [5:0] x3234_wVec_0_addr_0;
  wire [31:0] x3234_wVec_0_data;
  wire  x3234_wVec_0_en;
  wire  x3300_done;
  wire  x3300_en;
  wire  x3300_base_en;
  wire  x3300_mask;
  wire  x3300_resetter;
  wire  x3300_ctr_trivial;
  wire  x3238_valid_options_0;
  wire  x3238_valid_stops_0;
  wire  x3238_valid;
  wire [96:0] x3238_data_options_0;
  wire  x3238_ready;
  wire  x3240_ready_options_0;
  wire  x3240_ready;
  wire  x3240_now_valid;
  wire  x3240_valid;
  wire [31:0] x3240_0_number;
  wire  x3271_done;
  wire  x3271_en;
  wire  x3271_base_en;
  wire  x3271_mask;
  wire  x3271_resetter;
  wire  x3271_datapath_en;
  wire  x3271_ctr_trivial;
  wire [31:0] x3241_number;
  wire [31:0] x3242_number;
  wire [31:0] x3245_number;
  wire [31:0] x3246_number;
  wire [31:0] x3247_number;
  wire [31:0] x3248_number;
  wire [31:0] x3249_number;
  wire [31:0] x3252_number;
  wire  x3253;
  wire [31:0] x3254_number;
  wire [31:0] x3255_number;
  wire [31:0] x3256_number;
  wire [31:0] x3257_number;
  wire [31:0] x3258_number;
  wire [31:0] x3259_number;
  wire [31:0] x3260_number;
  wire [31:0] x3261_number;
  wire [31:0] x3262_number;
  wire [63:0] x3263_number;
  wire [63:0] x3265_number;
  wire [63:0] x3266_number;
  wire [63:0] x3267_item0;
  wire [31:0] x3267_item1;
  wire [96:0] x3267;
  wire [31:0] x3269_item0;
  wire [31:0] x3269_item1;
  wire [31:0] x3269_item2;
  wire [95:0] x3269;
  wire  x3299_done;
  wire  x3299_en;
  wire  x3299_base_en;
  wire  x3299_mask;
  wire  x3299_resetter;
  wire  x3299_ctr_trivial;
  wire  x3283_done;
  wire  x3283_en;
  wire  x3283_base_en;
  wire  x3283_mask;
  wire  x3283_resetter;
  wire  x3283_datapath_en;
  wire  x3283_ctr_trivial;
  wire [31:0] x3277_number;
  wire [31:0] x3279_number;
  wire [31:0] x3281_number;
  wire [31:0] x3284_number;
  wire  x3286_done;
  wire  x3286_en;
  wire  x3286_resetter;
  wire [31:0] x3285_0;
  wire  x3298_done;
  wire  x3298_en;
  wire  x3298_base_en;
  wire  x3298_mask;
  wire  x3298_datapath_en;
  wire  x3298_ctr_trivial;
  wire [31:0] b1331_number;
  wire [31:0] x3287_number;
  wire  x3288;
  wire [31:0] x3289_number;
  wire  x3290;
  wire  x3291;
  wire [31:0] x3292_number;
  wire  x3293;
  wire [31:0] x3295_number;
  wire  x3296;
  wire [5:0] x3297_wVec_0_addr_0;
  wire [31:0] x3297_wVec_0_data;
  wire  x3297_wVec_0_en;
  wire  x3428_done;
  wire  x3428_en;
  wire  x3428_base_en;
  wire  x3428_resetter;
  wire  x3428_ctr_trivial;
  wire  x3364_done;
  wire  x3364_en;
  wire  x3364_base_en;
  wire  x3364_mask;
  wire  x3364_resetter;
  wire  x3364_ctr_trivial;
  wire  x3302_valid_options_0;
  wire  x3302_valid_stops_0;
  wire  x3302_valid;
  wire [96:0] x3302_data_options_0;
  wire  x3302_ready;
  wire  x3304_ready_options_0;
  wire  x3304_ready;
  wire  x3304_now_valid;
  wire  x3304_valid;
  wire [31:0] x3304_0_number;
  wire  x3335_done;
  wire  x3335_en;
  wire  x3335_base_en;
  wire  x3335_mask;
  wire  x3335_resetter;
  wire  x3335_datapath_en;
  wire  x3335_ctr_trivial;
  wire [31:0] x3305_number;
  wire [31:0] x3306_number;
  wire [31:0] x3309_number;
  wire [31:0] x3310_number;
  wire [31:0] x3311_number;
  wire [31:0] x3312_number;
  wire [31:0] x3313_number;
  wire [31:0] x3316_number;
  wire  x3317;
  wire [31:0] x3318_number;
  wire [31:0] x3319_number;
  wire [31:0] x3320_number;
  wire [31:0] x3321_number;
  wire [31:0] x3322_number;
  wire [31:0] x3323_number;
  wire [31:0] x3324_number;
  wire [31:0] x3325_number;
  wire [31:0] x3326_number;
  wire [63:0] x3327_number;
  wire [63:0] x3329_number;
  wire [63:0] x3330_number;
  wire [63:0] x3331_item0;
  wire [31:0] x3331_item1;
  wire [96:0] x3331;
  wire [31:0] x3333_item0;
  wire [31:0] x3333_item1;
  wire [31:0] x3333_item2;
  wire [95:0] x3333;
  wire  x3363_done;
  wire  x3363_en;
  wire  x3363_base_en;
  wire  x3363_mask;
  wire  x3363_resetter;
  wire  x3363_ctr_trivial;
  wire  x3347_done;
  wire  x3347_en;
  wire  x3347_base_en;
  wire  x3347_mask;
  wire  x3347_resetter;
  wire  x3347_datapath_en;
  wire  x3347_ctr_trivial;
  wire [31:0] x3341_number;
  wire [31:0] x3343_number;
  wire [31:0] x3345_number;
  wire [31:0] x3348_number;
  wire  x3350_done;
  wire  x3350_en;
  wire  x3350_resetter;
  wire [31:0] x3349_0;
  wire  x3362_done;
  wire  x3362_en;
  wire  x3362_base_en;
  wire  x3362_mask;
  wire  x3362_datapath_en;
  wire  x3362_ctr_trivial;
  wire [31:0] b1393_number;
  wire [31:0] x3351_number;
  wire  x3352;
  wire [31:0] x3353_number;
  wire  x3354;
  wire  x3355;
  wire [31:0] x3356_number;
  wire  x3357;
  wire [31:0] x3359_number;
  wire  x3360;
  wire [5:0] x3361_wVec_0_addr_0;
  wire [31:0] x3361_wVec_0_data;
  wire  x3361_wVec_0_en;
  wire  x3427_done;
  wire  x3427_en;
  wire  x3427_base_en;
  wire  x3427_mask;
  wire  x3427_resetter;
  wire  x3427_ctr_trivial;
  wire  x3365_valid_options_0;
  wire  x3365_valid_stops_0;
  wire  x3365_valid;
  wire [96:0] x3365_data_options_0;
  wire  x3365_ready;
  wire  x3367_ready_options_0;
  wire  x3367_ready;
  wire  x3367_now_valid;
  wire  x3367_valid;
  wire [31:0] x3367_0_number;
  wire  x3398_done;
  wire  x3398_en;
  wire  x3398_base_en;
  wire  x3398_mask;
  wire  x3398_resetter;
  wire  x3398_datapath_en;
  wire  x3398_ctr_trivial;
  wire [31:0] x3368_number;
  wire [31:0] x3369_number;
  wire [31:0] x3372_number;
  wire [31:0] x3373_number;
  wire [31:0] x3374_number;
  wire [31:0] x3375_number;
  wire [31:0] x3376_number;
  wire [31:0] x3379_number;
  wire  x3380;
  wire [31:0] x3381_number;
  wire [31:0] x3382_number;
  wire [31:0] x3383_number;
  wire [31:0] x3384_number;
  wire [31:0] x3385_number;
  wire [31:0] x3386_number;
  wire [31:0] x3387_number;
  wire [31:0] x3388_number;
  wire [31:0] x3389_number;
  wire [63:0] x3390_number;
  wire [63:0] x3392_number;
  wire [63:0] x3393_number;
  wire [63:0] x3394_item0;
  wire [31:0] x3394_item1;
  wire [96:0] x3394;
  wire [31:0] x3396_item0;
  wire [31:0] x3396_item1;
  wire [31:0] x3396_item2;
  wire [95:0] x3396;
  wire  x3426_done;
  wire  x3426_en;
  wire  x3426_base_en;
  wire  x3426_mask;
  wire  x3426_resetter;
  wire  x3426_ctr_trivial;
  wire  x3410_done;
  wire  x3410_en;
  wire  x3410_base_en;
  wire  x3410_mask;
  wire  x3410_resetter;
  wire  x3410_datapath_en;
  wire  x3410_ctr_trivial;
  wire [31:0] x3404_number;
  wire [31:0] x3406_number;
  wire [31:0] x3408_number;
  wire [31:0] x3411_number;
  wire  x3413_done;
  wire  x3413_en;
  wire  x3413_resetter;
  wire [31:0] x3412_0;
  wire  x3425_done;
  wire  x3425_en;
  wire  x3425_base_en;
  wire  x3425_mask;
  wire  x3425_datapath_en;
  wire  x3425_ctr_trivial;
  wire [31:0] b1454_number;
  wire [31:0] x3414_number;
  wire  x3415;
  wire [31:0] x3416_number;
  wire  x3417;
  wire  x3418;
  wire [31:0] x3419_number;
  wire  x3420;
  wire [31:0] x3422_number;
  wire  x3423;
  wire [5:0] x3424_wVec_0_addr_0;
  wire [31:0] x3424_wVec_0_data;
  wire  x3424_wVec_0_en;
  wire  x3503_done;
  wire  x3503_en;
  wire  x3503_base_en;
  wire  x3503_resetter;
  wire  x3503_ctr_trivial;
  wire [31:0] x3431_number;
  wire  x3433_done;
  wire  x3433_en;
  wire  x3433_resetter;
  wire [31:0] x3432_0;
  wire [31:0] x3432_1;
  wire [31:0] x3432_2;
  wire [31:0] x3432_3;
  wire  x3466_done;
  wire  x3466_en;
  wire  x3466_base_en;
  wire  x3466_mask;
  wire  x3466_resetter;
  wire  x3466_datapath_en;
  wire  x3466_ctr_trivial;
  wire  x3466_rst_en;
  wire  x3429_wren;
  wire  x3429_resetter;
  wire [31:0] b1479_number;
  wire [31:0] b1480_number;
  wire [31:0] b1481_number;
  wire [31:0] b1482_number;
  wire  x3434;
  wire  x3435;
  wire  x3436;
  wire  x3437;
  wire [5:0] x3438_rVec_0_addr_0;
  wire  x3438_rVec_0_en;
  wire [5:0] x3438_rVec_1_addr_0;
  wire  x3438_rVec_1_en;
  wire [5:0] x3438_rVec_2_addr_0;
  wire  x3438_rVec_2_en;
  wire [5:0] x3438_rVec_3_addr_0;
  wire  x3438_rVec_3_en;
  wire [31:0] x3439_number;
  wire [31:0] x3440_number;
  wire [31:0] x3441_number;
  wire [31:0] x3442_number;
  wire [5:0] x3443_rVec_0_addr_0;
  wire  x3443_rVec_0_en;
  wire [5:0] x3443_rVec_1_addr_0;
  wire  x3443_rVec_1_en;
  wire [5:0] x3443_rVec_2_addr_0;
  wire  x3443_rVec_2_en;
  wire [5:0] x3443_rVec_3_addr_0;
  wire  x3443_rVec_3_en;
  wire [31:0] x3444_number;
  wire [31:0] x3445_number;
  wire [31:0] x3446_number;
  wire [31:0] x3447_number;
  wire [31:0] x3448_number;
  wire [31:0] x3449_number;
  wire [31:0] x3450_number;
  wire [31:0] x3451_number;
  wire [31:0] x3452_number;
  wire [31:0] x3453_number;
  wire [31:0] x3455_number;
  wire [31:0] x3456_number;
  wire  x3457;
  wire [31:0] x3458_number;
  wire [31:0] x3459_number;
  wire  x3462;
  wire [31:0] x3463_number;
  wire [31:0] x3464_number;
  wire [31:0] x3465_number;
  wire [31:0] x3467_number;
  wire  x3469_done;
  wire  x3469_en;
  wire  x3469_resetter;
  wire [31:0] x3468_0;
  wire [31:0] x3468_1;
  wire [31:0] x3468_2;
  wire [31:0] x3468_3;
  wire  x3502_done;
  wire  x3502_en;
  wire  x3502_base_en;
  wire  x3502_mask;
  wire  x3502_resetter;
  wire  x3502_datapath_en;
  wire  x3502_ctr_trivial;
  wire  x3502_rst_en;
  wire  x3430_wren;
  wire  x3430_resetter;
  wire [31:0] b1520_number;
  wire [31:0] b1521_number;
  wire [31:0] b1522_number;
  wire [31:0] b1523_number;
  wire  x3470;
  wire  x3471;
  wire  x3472;
  wire  x3473;
  wire [5:0] x3474_rVec_0_addr_0;
  wire  x3474_rVec_0_en;
  wire [5:0] x3474_rVec_1_addr_0;
  wire  x3474_rVec_1_en;
  wire [5:0] x3474_rVec_2_addr_0;
  wire  x3474_rVec_2_en;
  wire [5:0] x3474_rVec_3_addr_0;
  wire  x3474_rVec_3_en;
  wire [31:0] x3475_number;
  wire [31:0] x3476_number;
  wire [31:0] x3477_number;
  wire [31:0] x3478_number;
  wire [5:0] x3479_rVec_0_addr_0;
  wire  x3479_rVec_0_en;
  wire [5:0] x3479_rVec_1_addr_0;
  wire  x3479_rVec_1_en;
  wire [5:0] x3479_rVec_2_addr_0;
  wire  x3479_rVec_2_en;
  wire [5:0] x3479_rVec_3_addr_0;
  wire  x3479_rVec_3_en;
  wire [31:0] x3480_number;
  wire [31:0] x3481_number;
  wire [31:0] x3482_number;
  wire [31:0] x3483_number;
  wire [31:0] x3484_number;
  wire [31:0] x3485_number;
  wire [31:0] x3486_number;
  wire [31:0] x3487_number;
  wire [31:0] x3488_number;
  wire [31:0] x3489_number;
  wire [31:0] x3491_number;
  wire [31:0] x3492_number;
  wire  x3493;
  wire [31:0] x3494_number;
  wire [31:0] x3495_number;
  wire  x3498;
  wire [31:0] x3499_number;
  wire [31:0] x3500_number;
  wire [31:0] x3501_number;
  wire  x3514_done;
  wire  x3514_en;
  wire  x3514_base_en;
  wire  x3514_resetter;
  wire [31:0] x3504_number;
  wire [31:0] x3505_number;
  wire [31:0] x3506_number;
  wire [31:0] x3507_number;
  wire  x3510;
  wire [31:0] x3511_number;
  wire [31:0] x3512_number;
  wire [31:0] x3513_number;
  wire  x3518_done;
  wire  x3518_en;
  wire  x3518_base_en;
  wire  x3518_resetter;
  wire  x3518_datapath_en;
  wire  x3518_ctr_trivial;
  wire [31:0] x3516_number;
  wire  RootController_sm_clock;
  wire  RootController_sm_reset;
  wire  RootController_sm_io_input_enable;
  wire  RootController_sm_io_input_stageDone_0;
  wire  RootController_sm_io_input_stageDone_1;
  wire  RootController_sm_io_input_stageMask_0;
  wire  RootController_sm_io_input_stageMask_1;
  wire  RootController_sm_io_input_rst;
  wire  RootController_sm_io_output_done;
  wire  RootController_sm_io_output_stageEnable_0;
  wire  RootController_sm_io_output_stageEnable_1;
  wire  RootController_sm_io_output_rst_en;
  wire  x3152_0_clock;
  wire  x3152_0_reset;
  wire [31:0] x3152_0_io_input_0_data;
  wire [31:0] x3152_0_io_input_0_init;
  wire  x3152_0_io_input_0_enable;
  wire  x3152_0_io_input_0_reset;
  wire [31:0] x3152_0_io_output_data;
  wire  x3152_1_clock;
  wire  x3152_1_reset;
  wire [31:0] x3152_1_io_input_next;
  wire  x3152_1_io_input_enable;
  wire  x3152_1_io_input_reset;
  wire [31:0] x3152_1_io_output;
  wire  x3155_clock;
  wire  x3155_reset;
  wire [31:0] x3155_io_input_stops_0;
  wire  x3155_io_input_reset;
  wire  x3155_io_input_enable;
  wire [31:0] x3155_io_output_counts_1;
  wire [31:0] x3155_io_output_counts_0;
  wire  x3515_sm_clock;
  wire  x3515_sm_reset;
  wire  x3515_sm_io_input_enable;
  wire [31:0] x3515_sm_io_input_numIter;
  wire  x3515_sm_io_input_stageDone_0;
  wire  x3515_sm_io_input_stageDone_1;
  wire  x3515_sm_io_input_stageDone_2;
  wire  x3515_sm_io_input_stageDone_3;
  wire  x3515_sm_io_input_stageDone_4;
  wire  x3515_sm_io_input_rst;
  wire  x3515_sm_io_output_done;
  wire  x3515_sm_io_output_stageEnable_0;
  wire  x3515_sm_io_output_stageEnable_1;
  wire  x3515_sm_io_output_stageEnable_2;
  wire  x3515_sm_io_output_stageEnable_3;
  wire  x3515_sm_io_output_stageEnable_4;
  wire  x3515_sm_io_output_rst_en;
  wire  x3515_sm_io_output_ctr_inc;
  wire  b1204;
  wire  b1204_chain_read_1;
  wire  b1204_chain_read_2;
  wire  b1204_chain_read_3;
  wire  b1205;
  wire  b1205_chain_read_1;
  wire  b1205_chain_read_2;
  wire  b1205_chain_read_3;
  wire  b1205_chain_read_4;
  wire  b1202_chain_clock;
  wire  b1202_chain_reset;
  wire  b1202_chain_io_sEn_0;
  wire  b1202_chain_io_sEn_1;
  wire  b1202_chain_io_sEn_2;
  wire  b1202_chain_io_sEn_3;
  wire  b1202_chain_io_sEn_4;
  wire  b1202_chain_io_sDone_0;
  wire  b1202_chain_io_sDone_1;
  wire  b1202_chain_io_sDone_2;
  wire  b1202_chain_io_sDone_3;
  wire  b1202_chain_io_sDone_4;
  wire [31:0] b1202_chain_io_input_0_data;
  wire  b1202_chain_io_input_0_enable;
  wire  b1202_chain_io_input_0_reset;
  wire [31:0] b1202_chain_io_output_1_data;
  wire [31:0] b1202_chain_io_output_2_data;
  wire [31:0] b1202_chain_io_output_4_data;
  wire [31:0] b1202_chain_read_1;
  wire [31:0] b1202_chain_read_2;
  wire [31:0] b1202_chain_read_4;
  wire  b1203_chain_clock;
  wire  b1203_chain_reset;
  wire  b1203_chain_io_sEn_0;
  wire  b1203_chain_io_sEn_1;
  wire  b1203_chain_io_sEn_2;
  wire  b1203_chain_io_sEn_3;
  wire  b1203_chain_io_sEn_4;
  wire  b1203_chain_io_sDone_0;
  wire  b1203_chain_io_sDone_1;
  wire  b1203_chain_io_sDone_2;
  wire  b1203_chain_io_sDone_3;
  wire  b1203_chain_io_sDone_4;
  wire [31:0] b1203_chain_io_input_0_data;
  wire  b1203_chain_io_input_0_enable;
  wire  b1203_chain_io_input_0_reset;
  wire [31:0] b1203_chain_io_output_1_data;
  wire [31:0] b1203_chain_io_output_2_data;
  wire [31:0] b1203_chain_io_output_4_data;
  wire [31:0] b1203_chain_read_1;
  wire [31:0] b1203_chain_read_2;
  wire  x3156_0_clock;
  wire  x3156_0_reset;
  wire  x3156_0_io_sEn_0;
  wire  x3156_0_io_sEn_1;
  wire  x3156_0_io_sEn_2;
  wire  x3156_0_io_sEn_3;
  wire  x3156_0_io_sDone_0;
  wire  x3156_0_io_sDone_1;
  wire  x3156_0_io_sDone_2;
  wire  x3156_0_io_sDone_3;
  wire [31:0] x3156_0_io_input_0_data;
  wire  x3156_0_io_input_0_enable;
  wire  x3156_0_io_input_0_reset;
  wire [31:0] x3156_0_io_output_1_data;
  wire [31:0] x3156_0_io_output_2_data;
  wire [31:0] x3156_0_io_output_3_data;
  wire  x3157_0_clock;
  wire  x3157_0_reset;
  wire  x3157_0_io_sEn_0;
  wire  x3157_0_io_sEn_1;
  wire  x3157_0_io_sEn_2;
  wire  x3157_0_io_sEn_3;
  wire  x3157_0_io_sDone_0;
  wire  x3157_0_io_sDone_1;
  wire  x3157_0_io_sDone_2;
  wire  x3157_0_io_sDone_3;
  wire [31:0] x3157_0_io_input_0_data;
  wire  x3157_0_io_input_0_enable;
  wire  x3157_0_io_input_0_reset;
  wire [31:0] x3157_0_io_output_1_data;
  wire [31:0] x3157_0_io_output_2_data;
  wire [31:0] x3157_0_io_output_3_data;
  wire  x3158_0_clock;
  wire  x3158_0_reset;
  wire  x3158_0_io_sEn_0;
  wire  x3158_0_io_sEn_1;
  wire  x3158_0_io_sEn_2;
  wire  x3158_0_io_sDone_0;
  wire  x3158_0_io_sDone_1;
  wire  x3158_0_io_sDone_2;
  wire [5:0] x3158_0_io_w_0_addr_0;
  wire [31:0] x3158_0_io_w_0_data;
  wire  x3158_0_io_w_0_en;
  wire [5:0] x3158_0_io_r_0_addr_0;
  wire  x3158_0_io_r_0_en;
  wire [5:0] x3158_0_io_r_1_addr_0;
  wire  x3158_0_io_r_1_en;
  wire [5:0] x3158_0_io_r_2_addr_0;
  wire  x3158_0_io_r_2_en;
  wire [5:0] x3158_0_io_r_3_addr_0;
  wire  x3158_0_io_r_3_en;
  wire [31:0] x3158_0_io_output_data_8;
  wire [31:0] x3158_0_io_output_data_9;
  wire [31:0] x3158_0_io_output_data_10;
  wire [31:0] x3158_0_io_output_data_11;
  wire  x3159_0_clock;
  wire  x3159_0_reset;
  wire  x3159_0_io_sEn_0;
  wire  x3159_0_io_sEn_1;
  wire  x3159_0_io_sEn_2;
  wire  x3159_0_io_sDone_0;
  wire  x3159_0_io_sDone_1;
  wire  x3159_0_io_sDone_2;
  wire [5:0] x3159_0_io_w_0_addr_0;
  wire [31:0] x3159_0_io_w_0_data;
  wire  x3159_0_io_w_0_en;
  wire [5:0] x3159_0_io_r_0_addr_0;
  wire  x3159_0_io_r_0_en;
  wire [5:0] x3159_0_io_r_1_addr_0;
  wire  x3159_0_io_r_1_en;
  wire [5:0] x3159_0_io_r_2_addr_0;
  wire  x3159_0_io_r_2_en;
  wire [5:0] x3159_0_io_r_3_addr_0;
  wire  x3159_0_io_r_3_en;
  wire [31:0] x3159_0_io_output_data_8;
  wire [31:0] x3159_0_io_output_data_9;
  wire [31:0] x3159_0_io_output_data_10;
  wire [31:0] x3159_0_io_output_data_11;
  wire  x3160_0_clock;
  wire  x3160_0_reset;
  wire  x3160_0_io_sEn_0;
  wire  x3160_0_io_sEn_1;
  wire  x3160_0_io_sDone_0;
  wire  x3160_0_io_sDone_1;
  wire [5:0] x3160_0_io_w_0_addr_0;
  wire [31:0] x3160_0_io_w_0_data;
  wire  x3160_0_io_w_0_en;
  wire [5:0] x3160_0_io_r_0_addr_0;
  wire  x3160_0_io_r_0_en;
  wire [5:0] x3160_0_io_r_1_addr_0;
  wire  x3160_0_io_r_1_en;
  wire [5:0] x3160_0_io_r_2_addr_0;
  wire  x3160_0_io_r_2_en;
  wire [5:0] x3160_0_io_r_3_addr_0;
  wire  x3160_0_io_r_3_en;
  wire [31:0] x3160_0_io_output_data_4;
  wire [31:0] x3160_0_io_output_data_5;
  wire [31:0] x3160_0_io_output_data_6;
  wire [31:0] x3160_0_io_output_data_7;
  wire  x3161_0_clock;
  wire  x3161_0_reset;
  wire  x3161_0_io_sEn_0;
  wire  x3161_0_io_sEn_1;
  wire  x3161_0_io_sDone_0;
  wire  x3161_0_io_sDone_1;
  wire [5:0] x3161_0_io_w_0_addr_0;
  wire [31:0] x3161_0_io_w_0_data;
  wire  x3161_0_io_w_0_en;
  wire [5:0] x3161_0_io_r_0_addr_0;
  wire  x3161_0_io_r_0_en;
  wire [5:0] x3161_0_io_r_1_addr_0;
  wire  x3161_0_io_r_1_en;
  wire [5:0] x3161_0_io_r_2_addr_0;
  wire  x3161_0_io_r_2_en;
  wire [5:0] x3161_0_io_r_3_addr_0;
  wire  x3161_0_io_r_3_en;
  wire [31:0] x3161_0_io_output_data_4;
  wire [31:0] x3161_0_io_output_data_5;
  wire [31:0] x3161_0_io_output_data_6;
  wire [31:0] x3161_0_io_output_data_7;
  wire  x3174_sm_clock;
  wire  x3174_sm_reset;
  wire  x3174_sm_io_input_enable;
  wire  x3174_sm_io_input_stageDone_0;
  wire  x3174_sm_io_input_stageDone_1;
  wire  x3174_sm_io_input_stageMask_0;
  wire  x3174_sm_io_input_stageMask_1;
  wire  x3174_sm_io_input_rst;
  wire  x3174_sm_io_output_done;
  wire  x3174_sm_io_output_stageEnable_0;
  wire  x3174_sm_io_output_stageEnable_1;
  wire  x3174_sm_io_output_rst_en;
  wire  x3167_sm_clock;
  wire  x3167_sm_reset;
  wire  x3167_sm_io_input_enable;
  wire  x3167_sm_io_input_ctr_done;
  wire  x3167_sm_io_input_rst;
  wire  x3167_sm_io_output_done;
  wire  x3167_sm_io_output_ctr_inc;
  wire  x3173_sm_clock;
  wire  x3173_sm_reset;
  wire  x3173_sm_io_input_enable;
  wire  x3173_sm_io_input_ctr_done;
  wire  x3173_sm_io_input_rst;
  wire  x3173_sm_io_output_done;
  wire  x3173_sm_io_output_ctr_inc;
  wire  x3301_sm_clock;
  wire  x3301_sm_reset;
  wire  x3301_sm_io_input_enable;
  wire  x3301_sm_io_input_stageDone_0;
  wire  x3301_sm_io_input_stageDone_1;
  wire  x3301_sm_io_input_stageMask_0;
  wire  x3301_sm_io_input_stageMask_1;
  wire  x3301_sm_io_input_rst;
  wire  x3301_sm_io_output_done;
  wire  x3301_sm_io_output_stageEnable_0;
  wire  x3301_sm_io_output_stageEnable_1;
  wire  x3301_sm_io_output_rst_en;
  wire  x3237_sm_clock;
  wire  x3237_sm_reset;
  wire  x3237_sm_io_input_enable;
  wire  x3237_sm_io_input_stageDone_0;
  wire  x3237_sm_io_input_stageDone_1;
  wire  x3237_sm_io_input_stageMask_0;
  wire  x3237_sm_io_input_stageMask_1;
  wire  x3237_sm_io_input_rst;
  wire  x3237_sm_io_output_done;
  wire  x3237_sm_io_output_stageEnable_0;
  wire  x3237_sm_io_output_stageEnable_1;
  wire  x3237_sm_io_output_rst_en;
  wire  x3175_valid_srff_clock;
  wire  x3175_valid_srff_reset;
  wire  x3175_valid_srff_io_input_set;
  wire  x3175_valid_srff_io_input_reset;
  wire  x3175_valid_srff_io_input_asyn_reset;
  wire  x3175_valid_srff_io_output_data;
  wire  _T_1601;
  wire  x3176_clock;
  wire  x3176_reset;
  wire [95:0] x3176_io_in_0_data;
  wire  x3176_io_in_0_en;
  wire [95:0] x3176_io_out_0;
  wire  x3176_io_deq_0;
  wire  x3176_io_empty;
  wire  x3176_io_full;
  wire  x3208_sm_clock;
  wire  x3208_sm_reset;
  wire  x3208_sm_io_input_enable;
  wire  x3208_sm_io_input_ctr_done;
  wire  x3208_sm_io_input_rst;
  wire  x3208_sm_io_output_done;
  wire  x3208_sm_io_output_ctr_inc;
  wire  x3236_sm_clock;
  wire  x3236_sm_reset;
  wire  x3236_sm_io_input_enable;
  wire  x3236_sm_io_input_stageDone_0;
  wire  x3236_sm_io_input_stageDone_1;
  wire  x3236_sm_io_input_stageMask_0;
  wire  x3236_sm_io_input_stageMask_1;
  wire  x3236_sm_io_input_rst;
  wire  x3236_sm_io_output_done;
  wire  x3236_sm_io_output_stageEnable_0;
  wire  x3236_sm_io_output_stageEnable_1;
  wire  x3236_sm_io_output_rst_en;
  wire  x3210_0_clock;
  wire  x3210_0_reset;
  wire [31:0] x3210_0_io_input_0_data;
  wire [31:0] x3210_0_io_input_0_init;
  wire  x3210_0_io_input_0_enable;
  wire  x3210_0_io_input_0_reset;
  wire [31:0] x3210_0_io_output_data;
  wire  x3211_0_clock;
  wire  x3211_0_reset;
  wire [31:0] x3211_0_io_input_0_data;
  wire [31:0] x3211_0_io_input_0_init;
  wire  x3211_0_io_input_0_enable;
  wire  x3211_0_io_input_0_reset;
  wire [31:0] x3211_0_io_output_data;
  wire  x3212_0_clock;
  wire  x3212_0_reset;
  wire [31:0] x3212_0_io_input_0_data;
  wire [31:0] x3212_0_io_input_0_init;
  wire  x3212_0_io_input_0_enable;
  wire  x3212_0_io_input_0_reset;
  wire [31:0] x3212_0_io_output_data;
  wire  x3220_sm_clock;
  wire  x3220_sm_reset;
  wire  x3220_sm_io_input_enable;
  wire  x3220_sm_io_input_ctr_done;
  wire  x3220_sm_io_input_rst;
  wire  x3220_sm_io_output_done;
  wire  x3220_sm_io_output_ctr_inc;
  wire  x3223_clock;
  wire  x3223_reset;
  wire [31:0] x3223_io_input_stops_0;
  wire  x3223_io_input_reset;
  wire  x3223_io_input_enable;
  wire [31:0] x3223_io_output_counts_0;
  wire  x3223_io_output_done;
  wire  x3235_sm_io_input_ctr_done;
  wire  x3235_sm_io_output_done;
  wire  b1271;
  wire  x3300_sm_clock;
  wire  x3300_sm_reset;
  wire  x3300_sm_io_input_enable;
  wire  x3300_sm_io_input_stageDone_0;
  wire  x3300_sm_io_input_stageDone_1;
  wire  x3300_sm_io_input_stageMask_0;
  wire  x3300_sm_io_input_stageMask_1;
  wire  x3300_sm_io_input_rst;
  wire  x3300_sm_io_output_done;
  wire  x3300_sm_io_output_stageEnable_0;
  wire  x3300_sm_io_output_stageEnable_1;
  wire  x3300_sm_io_output_rst_en;
  wire  x3238_valid_srff_clock;
  wire  x3238_valid_srff_reset;
  wire  x3238_valid_srff_io_input_set;
  wire  x3238_valid_srff_io_input_reset;
  wire  x3238_valid_srff_io_input_asyn_reset;
  wire  x3238_valid_srff_io_output_data;
  wire  _T_1610;
  wire  x3239_clock;
  wire  x3239_reset;
  wire [95:0] x3239_io_in_0_data;
  wire  x3239_io_in_0_en;
  wire [95:0] x3239_io_out_0;
  wire  x3239_io_deq_0;
  wire  x3239_io_empty;
  wire  x3239_io_full;
  wire  x3271_sm_clock;
  wire  x3271_sm_reset;
  wire  x3271_sm_io_input_enable;
  wire  x3271_sm_io_input_ctr_done;
  wire  x3271_sm_io_input_rst;
  wire  x3271_sm_io_output_done;
  wire  x3271_sm_io_output_ctr_inc;
  wire  x3299_sm_clock;
  wire  x3299_sm_reset;
  wire  x3299_sm_io_input_enable;
  wire  x3299_sm_io_input_stageDone_0;
  wire  x3299_sm_io_input_stageDone_1;
  wire  x3299_sm_io_input_stageMask_0;
  wire  x3299_sm_io_input_stageMask_1;
  wire  x3299_sm_io_input_rst;
  wire  x3299_sm_io_output_done;
  wire  x3299_sm_io_output_stageEnable_0;
  wire  x3299_sm_io_output_stageEnable_1;
  wire  x3299_sm_io_output_rst_en;
  wire  x3273_0_clock;
  wire  x3273_0_reset;
  wire [31:0] x3273_0_io_input_0_data;
  wire [31:0] x3273_0_io_input_0_init;
  wire  x3273_0_io_input_0_enable;
  wire  x3273_0_io_input_0_reset;
  wire [31:0] x3273_0_io_output_data;
  wire  x3274_0_clock;
  wire  x3274_0_reset;
  wire [31:0] x3274_0_io_input_0_data;
  wire [31:0] x3274_0_io_input_0_init;
  wire  x3274_0_io_input_0_enable;
  wire  x3274_0_io_input_0_reset;
  wire [31:0] x3274_0_io_output_data;
  wire  x3275_0_clock;
  wire  x3275_0_reset;
  wire [31:0] x3275_0_io_input_0_data;
  wire [31:0] x3275_0_io_input_0_init;
  wire  x3275_0_io_input_0_enable;
  wire  x3275_0_io_input_0_reset;
  wire [31:0] x3275_0_io_output_data;
  wire  x3283_sm_clock;
  wire  x3283_sm_reset;
  wire  x3283_sm_io_input_enable;
  wire  x3283_sm_io_input_ctr_done;
  wire  x3283_sm_io_input_rst;
  wire  x3283_sm_io_output_done;
  wire  x3283_sm_io_output_ctr_inc;
  wire  x3286_clock;
  wire  x3286_reset;
  wire [31:0] x3286_io_input_stops_0;
  wire  x3286_io_input_reset;
  wire  x3286_io_input_enable;
  wire [31:0] x3286_io_output_counts_0;
  wire  x3286_io_output_done;
  wire  x3298_sm_io_input_ctr_done;
  wire  x3298_sm_io_output_done;
  wire  b1332;
  wire  x3428_sm_clock;
  wire  x3428_sm_reset;
  wire  x3428_sm_io_input_enable;
  wire  x3428_sm_io_input_stageDone_0;
  wire  x3428_sm_io_input_stageDone_1;
  wire  x3428_sm_io_input_stageMask_0;
  wire  x3428_sm_io_input_stageMask_1;
  wire  x3428_sm_io_input_rst;
  wire  x3428_sm_io_output_done;
  wire  x3428_sm_io_output_stageEnable_0;
  wire  x3428_sm_io_output_stageEnable_1;
  wire  x3428_sm_io_output_rst_en;
  wire  x3364_sm_clock;
  wire  x3364_sm_reset;
  wire  x3364_sm_io_input_enable;
  wire  x3364_sm_io_input_stageDone_0;
  wire  x3364_sm_io_input_stageDone_1;
  wire  x3364_sm_io_input_stageMask_0;
  wire  x3364_sm_io_input_stageMask_1;
  wire  x3364_sm_io_input_rst;
  wire  x3364_sm_io_output_done;
  wire  x3364_sm_io_output_stageEnable_0;
  wire  x3364_sm_io_output_stageEnable_1;
  wire  x3364_sm_io_output_rst_en;
  wire  x3302_valid_srff_clock;
  wire  x3302_valid_srff_reset;
  wire  x3302_valid_srff_io_input_set;
  wire  x3302_valid_srff_io_input_reset;
  wire  x3302_valid_srff_io_input_asyn_reset;
  wire  x3302_valid_srff_io_output_data;
  wire  _T_1619;
  wire  x3303_clock;
  wire  x3303_reset;
  wire [95:0] x3303_io_in_0_data;
  wire  x3303_io_in_0_en;
  wire [95:0] x3303_io_out_0;
  wire  x3303_io_deq_0;
  wire  x3303_io_empty;
  wire  x3303_io_full;
  wire  x3335_sm_clock;
  wire  x3335_sm_reset;
  wire  x3335_sm_io_input_enable;
  wire  x3335_sm_io_input_ctr_done;
  wire  x3335_sm_io_input_rst;
  wire  x3335_sm_io_output_done;
  wire  x3335_sm_io_output_ctr_inc;
  wire  x3363_sm_clock;
  wire  x3363_sm_reset;
  wire  x3363_sm_io_input_enable;
  wire  x3363_sm_io_input_stageDone_0;
  wire  x3363_sm_io_input_stageDone_1;
  wire  x3363_sm_io_input_stageMask_0;
  wire  x3363_sm_io_input_stageMask_1;
  wire  x3363_sm_io_input_rst;
  wire  x3363_sm_io_output_done;
  wire  x3363_sm_io_output_stageEnable_0;
  wire  x3363_sm_io_output_stageEnable_1;
  wire  x3363_sm_io_output_rst_en;
  wire  x3337_0_clock;
  wire  x3337_0_reset;
  wire [31:0] x3337_0_io_input_0_data;
  wire [31:0] x3337_0_io_input_0_init;
  wire  x3337_0_io_input_0_enable;
  wire  x3337_0_io_input_0_reset;
  wire [31:0] x3337_0_io_output_data;
  wire  x3338_0_clock;
  wire  x3338_0_reset;
  wire [31:0] x3338_0_io_input_0_data;
  wire [31:0] x3338_0_io_input_0_init;
  wire  x3338_0_io_input_0_enable;
  wire  x3338_0_io_input_0_reset;
  wire [31:0] x3338_0_io_output_data;
  wire  x3339_0_clock;
  wire  x3339_0_reset;
  wire [31:0] x3339_0_io_input_0_data;
  wire [31:0] x3339_0_io_input_0_init;
  wire  x3339_0_io_input_0_enable;
  wire  x3339_0_io_input_0_reset;
  wire [31:0] x3339_0_io_output_data;
  wire  x3347_sm_clock;
  wire  x3347_sm_reset;
  wire  x3347_sm_io_input_enable;
  wire  x3347_sm_io_input_ctr_done;
  wire  x3347_sm_io_input_rst;
  wire  x3347_sm_io_output_done;
  wire  x3347_sm_io_output_ctr_inc;
  wire  x3350_clock;
  wire  x3350_reset;
  wire [31:0] x3350_io_input_stops_0;
  wire  x3350_io_input_reset;
  wire  x3350_io_input_enable;
  wire [31:0] x3350_io_output_counts_0;
  wire  x3350_io_output_done;
  wire  x3362_sm_io_input_ctr_done;
  wire  x3362_sm_io_output_done;
  wire  b1394;
  wire  x3427_sm_clock;
  wire  x3427_sm_reset;
  wire  x3427_sm_io_input_enable;
  wire  x3427_sm_io_input_stageDone_0;
  wire  x3427_sm_io_input_stageDone_1;
  wire  x3427_sm_io_input_stageMask_0;
  wire  x3427_sm_io_input_stageMask_1;
  wire  x3427_sm_io_input_rst;
  wire  x3427_sm_io_output_done;
  wire  x3427_sm_io_output_stageEnable_0;
  wire  x3427_sm_io_output_stageEnable_1;
  wire  x3427_sm_io_output_rst_en;
  wire  x3365_valid_srff_clock;
  wire  x3365_valid_srff_reset;
  wire  x3365_valid_srff_io_input_set;
  wire  x3365_valid_srff_io_input_reset;
  wire  x3365_valid_srff_io_input_asyn_reset;
  wire  x3365_valid_srff_io_output_data;
  wire  _T_1628;
  wire  x3366_clock;
  wire  x3366_reset;
  wire [95:0] x3366_io_in_0_data;
  wire  x3366_io_in_0_en;
  wire [95:0] x3366_io_out_0;
  wire  x3366_io_deq_0;
  wire  x3366_io_empty;
  wire  x3366_io_full;
  wire  x3398_sm_clock;
  wire  x3398_sm_reset;
  wire  x3398_sm_io_input_enable;
  wire  x3398_sm_io_input_ctr_done;
  wire  x3398_sm_io_input_rst;
  wire  x3398_sm_io_output_done;
  wire  x3398_sm_io_output_ctr_inc;
  wire  x3426_sm_clock;
  wire  x3426_sm_reset;
  wire  x3426_sm_io_input_enable;
  wire  x3426_sm_io_input_stageDone_0;
  wire  x3426_sm_io_input_stageDone_1;
  wire  x3426_sm_io_input_stageMask_0;
  wire  x3426_sm_io_input_stageMask_1;
  wire  x3426_sm_io_input_rst;
  wire  x3426_sm_io_output_done;
  wire  x3426_sm_io_output_stageEnable_0;
  wire  x3426_sm_io_output_stageEnable_1;
  wire  x3426_sm_io_output_rst_en;
  wire  x3400_0_clock;
  wire  x3400_0_reset;
  wire [31:0] x3400_0_io_input_0_data;
  wire [31:0] x3400_0_io_input_0_init;
  wire  x3400_0_io_input_0_enable;
  wire  x3400_0_io_input_0_reset;
  wire [31:0] x3400_0_io_output_data;
  wire  x3401_0_clock;
  wire  x3401_0_reset;
  wire [31:0] x3401_0_io_input_0_data;
  wire [31:0] x3401_0_io_input_0_init;
  wire  x3401_0_io_input_0_enable;
  wire  x3401_0_io_input_0_reset;
  wire [31:0] x3401_0_io_output_data;
  wire  x3402_0_clock;
  wire  x3402_0_reset;
  wire [31:0] x3402_0_io_input_0_data;
  wire [31:0] x3402_0_io_input_0_init;
  wire  x3402_0_io_input_0_enable;
  wire  x3402_0_io_input_0_reset;
  wire [31:0] x3402_0_io_output_data;
  wire  x3410_sm_clock;
  wire  x3410_sm_reset;
  wire  x3410_sm_io_input_enable;
  wire  x3410_sm_io_input_ctr_done;
  wire  x3410_sm_io_input_rst;
  wire  x3410_sm_io_output_done;
  wire  x3410_sm_io_output_ctr_inc;
  wire  x3413_clock;
  wire  x3413_reset;
  wire [31:0] x3413_io_input_stops_0;
  wire  x3413_io_input_reset;
  wire  x3413_io_input_enable;
  wire [31:0] x3413_io_output_counts_0;
  wire  x3413_io_output_done;
  wire  x3425_sm_io_input_ctr_done;
  wire  x3425_sm_io_output_done;
  wire  b1455;
  wire  x3429_0_clock;
  wire  x3429_0_reset;
  wire [31:0] x3429_0_io_input_next;
  wire  x3429_0_io_input_enable;
  wire  x3429_0_io_input_reset;
  wire [31:0] x3429_0_io_output;
  wire  x3429_1_clock;
  wire  x3429_1_reset;
  wire  x3429_1_io_sEn_0;
  wire  x3429_1_io_sEn_1;
  wire  x3429_1_io_sDone_0;
  wire  x3429_1_io_sDone_1;
  wire [31:0] x3429_1_io_input_0_data;
  wire  x3429_1_io_input_0_enable;
  wire  x3429_1_io_input_0_reset;
  wire [31:0] x3429_1_io_output_1_data;
  wire  x3430_0_clock;
  wire  x3430_0_reset;
  wire [31:0] x3430_0_io_input_next;
  wire  x3430_0_io_input_enable;
  wire  x3430_0_io_input_reset;
  wire [31:0] x3430_0_io_output;
  wire  x3430_1_clock;
  wire  x3430_1_reset;
  wire  x3430_1_io_sEn_0;
  wire  x3430_1_io_sEn_1;
  wire  x3430_1_io_sDone_0;
  wire  x3430_1_io_sDone_1;
  wire [31:0] x3430_1_io_input_0_data;
  wire  x3430_1_io_input_0_enable;
  wire  x3430_1_io_input_0_reset;
  wire [31:0] x3430_1_io_output_1_data;
  wire  x3503_sm_clock;
  wire  x3503_sm_reset;
  wire  x3503_sm_io_input_enable;
  wire  x3503_sm_io_input_stageDone_0;
  wire  x3503_sm_io_input_stageDone_1;
  wire  x3503_sm_io_input_stageMask_0;
  wire  x3503_sm_io_input_stageMask_1;
  wire  x3503_sm_io_input_rst;
  wire  x3503_sm_io_output_done;
  wire  x3503_sm_io_output_stageEnable_0;
  wire  x3503_sm_io_output_stageEnable_1;
  wire  x3503_sm_io_output_rst_en;
  wire  x3433_clock;
  wire  x3433_reset;
  wire [31:0] x3433_io_input_stops_0;
  wire  x3433_io_input_reset;
  wire  x3433_io_input_enable;
  wire [31:0] x3433_io_output_counts_3;
  wire [31:0] x3433_io_output_counts_2;
  wire [31:0] x3433_io_output_counts_1;
  wire [31:0] x3433_io_output_counts_0;
  wire  x3433_io_output_done;
  wire  x3466_sm_clock;
  wire  x3466_sm_reset;
  wire  x3466_sm_io_input_enable;
  wire  x3466_sm_io_input_ctr_done;
  wire  x3466_sm_io_input_rst;
  wire  x3466_sm_io_output_done;
  wire  x3466_sm_io_output_ctr_inc;
  wire  x3466_sm_io_output_rst_en;
  wire  b1483;
  wire  b1484;
  wire  b1485;
  wire  b1486;
  wire  x3469_clock;
  wire  x3469_reset;
  wire [31:0] x3469_io_input_stops_0;
  wire  x3469_io_input_reset;
  wire  x3469_io_input_enable;
  wire [31:0] x3469_io_output_counts_3;
  wire [31:0] x3469_io_output_counts_2;
  wire [31:0] x3469_io_output_counts_1;
  wire [31:0] x3469_io_output_counts_0;
  wire  x3469_io_output_done;
  wire  x3502_sm_clock;
  wire  x3502_sm_reset;
  wire  x3502_sm_io_input_enable;
  wire  x3502_sm_io_input_ctr_done;
  wire  x3502_sm_io_input_rst;
  wire  x3502_sm_io_output_done;
  wire  x3502_sm_io_output_ctr_inc;
  wire  x3502_sm_io_output_rst_en;
  wire  b1524;
  wire  b1525;
  wire  b1526;
  wire  b1527;
  wire  x3514_sm_clock;
  wire  x3514_sm_reset;
  wire  x3514_sm_io_input_enable;
  wire  x3514_sm_io_input_ctr_done;
  wire  x3514_sm_io_input_rst;
  wire  x3514_sm_io_output_done;
  wire  x3514_sm_io_output_ctr_inc;
  wire  b1204_chain_clock;
  wire  b1204_chain_reset;
  wire  b1204_chain_io_sEn_0;
  wire  b1204_chain_io_sEn_1;
  wire  b1204_chain_io_sEn_2;
  wire  b1204_chain_io_sEn_3;
  wire  b1204_chain_io_sEn_4;
  wire  b1204_chain_io_sDone_0;
  wire  b1204_chain_io_sDone_1;
  wire  b1204_chain_io_sDone_2;
  wire  b1204_chain_io_sDone_3;
  wire  b1204_chain_io_sDone_4;
  wire  b1204_chain_io_input_0_data;
  wire  b1204_chain_io_input_0_enable;
  wire  b1204_chain_io_input_0_reset;
  wire  b1204_chain_io_output_1_data;
  wire  b1204_chain_io_output_2_data;
  wire  b1204_chain_io_output_3_data;
  wire  b1204_chain_io_output_4_data;
  wire  _T_1660;
  wire  _T_1662;
  wire  _T_1664;
  wire  b1205_chain_clock;
  wire  b1205_chain_reset;
  wire  b1205_chain_io_sEn_0;
  wire  b1205_chain_io_sEn_1;
  wire  b1205_chain_io_sEn_2;
  wire  b1205_chain_io_sEn_3;
  wire  b1205_chain_io_sEn_4;
  wire  b1205_chain_io_sDone_0;
  wire  b1205_chain_io_sDone_1;
  wire  b1205_chain_io_sDone_2;
  wire  b1205_chain_io_sDone_3;
  wire  b1205_chain_io_sDone_4;
  wire  b1205_chain_io_input_0_data;
  wire  b1205_chain_io_input_0_enable;
  wire  b1205_chain_io_input_0_reset;
  wire  b1205_chain_io_output_1_data;
  wire  b1205_chain_io_output_2_data;
  wire  b1205_chain_io_output_3_data;
  wire  b1205_chain_io_output_4_data;
  wire  _T_1668;
  wire  _T_1670;
  wire  _T_1672;
  wire  _T_1674;
  wire  x3518_sm_clock;
  wire  x3518_sm_reset;
  wire  x3518_sm_io_input_enable;
  wire  x3518_sm_io_input_ctr_done;
  wire  x3518_sm_io_input_rst;
  wire  x3518_sm_io_output_done;
  wire  x3518_sm_io_output_ctr_inc;
  wire  _T_1675;
  wire  _T_1678;
  wire  _T_1679;
  reg  _T_1682;
  reg [31:0] _RAND_0;
  wire  _T_1688;
  wire  _T_1697;
  wire  _T_1698;
  wire  RetimeWrapper_1_clock;
  wire  RetimeWrapper_1_reset;
  wire  RetimeWrapper_1_io_flow;
  wire  RetimeWrapper_1_io_in;
  wire  RetimeWrapper_1_io_out;
  wire  _T_1702;
  wire  retime_counter_clock;
  wire  retime_counter_reset;
  wire  retime_counter_io_input_reset;
  wire  retime_counter_io_output_done;
  wire  RetimeWrapper_2_clock;
  wire  RetimeWrapper_2_reset;
  wire  RetimeWrapper_2_io_flow;
  wire  RetimeWrapper_2_io_in;
  wire  RetimeWrapper_2_io_out;
  wire  _T_1710;
  wire [31:0] _T_1711;
  wire [32:0] _T_1722_number;
  wire [32:0] _T_1724_number;
  wire [32:0] _T_1734;
  wire  _T_1737;
  wire [32:0] _T_1739;
  wire [33:0] _T_1753;
  wire [33:0] _T_1754;
  wire [32:0] _T_1755;
  wire [31:0] x35150_range_number;
  wire [31:0] _T_1770;
  wire [31:0] _T_1774;
  wire [31:0] _T_1780;
  wire [32:0] _T_1782;
  wire [31:0] x35150_hops_number;
  wire [32:0] _T_1784;
  wire [31:0] _T_1786_number;
  wire [31:0] _T_1788_number;
  wire [31:0] _T_1796;
  wire [63:0] _T_1805_number;
  wire [31:0] _GEN_8;
  wire [31:0] _T_1806;
  wire [31:0] x35150_leftover_number;
  wire [31:0] _T_1815;
  wire [31:0] _T_1881;
  wire  x35150_evenfit;
  wire  x35150_adjustment;
  wire [31:0] _T_1909_number;
  wire  _T_1911_number;
  wire [31:0] _T_1919;
  wire [31:0] _T_1928;
  wire [32:0] _T_1930_number;
  wire [32:0] _T_1932_number;
  wire [32:0] _T_1934_number;
  wire [32:0] _T_1942;
  wire [32:0] _T_1947;
  wire [32:0] _T_1955;
  wire [32:0] _T_1960;
  wire [33:0] _T_1961;
  wire [32:0] _T_1962;
  wire [31:0] _T_1964_number;
  wire [31:0] _T_1972;
  wire [31:0] _T_1976;
  wire  _T_1978;
  wire  _T_1981;
  wire  _T_1982;
  reg  _T_1985;
  reg [31:0] _RAND_1;
  wire  _T_1991;
  wire  _T_1992;
  wire  _T_1996;
  wire  _T_1999;
  wire [31:0] _T_2075_number;
  wire [31:0] _T_2077_number;
  wire [31:0] _T_2085;
  wire [31:0] _T_2096;
  wire [31:0] _T_2100;
  wire [31:0] _T_2101;
  wire  _T_2102;
  wire  RetimeWrapper_3_clock;
  wire  RetimeWrapper_3_reset;
  wire  RetimeWrapper_3_io_flow;
  wire  RetimeWrapper_3_io_in;
  wire  RetimeWrapper_3_io_out;
  wire  _T_2136;
  wire [31:0] _T_2212_number;
  wire [31:0] _T_2214_number;
  wire [31:0] _T_2222;
  wire [31:0] _T_2233;
  wire [31:0] _T_2237;
  wire [31:0] _T_2238;
  wire  _T_2239;
  wire  RetimeWrapper_4_clock;
  wire  RetimeWrapper_4_reset;
  wire  RetimeWrapper_4_io_flow;
  wire  RetimeWrapper_4_io_in;
  wire  RetimeWrapper_4_io_out;
  wire  _T_2273;
  wire  RetimeWrapper_5_clock;
  wire  RetimeWrapper_5_reset;
  wire  RetimeWrapper_5_io_flow;
  wire  RetimeWrapper_5_io_in;
  wire  RetimeWrapper_5_io_out;
  wire  _T_2280;
  wire  _T_2282;
  wire  _T_2283;
  wire  RetimeWrapper_6_clock;
  wire  RetimeWrapper_6_reset;
  wire  RetimeWrapper_6_io_flow;
  wire  RetimeWrapper_6_io_in;
  wire  RetimeWrapper_6_io_out;
  wire  _T_2287;
  wire  _T_2289;
  wire  _T_2290;
  wire  RetimeWrapper_7_clock;
  wire  RetimeWrapper_7_reset;
  wire  RetimeWrapper_7_io_flow;
  wire  RetimeWrapper_7_io_in;
  wire  RetimeWrapper_7_io_out;
  wire  _T_2294;
  wire  _T_2296;
  wire  RetimeWrapper_8_clock;
  wire  RetimeWrapper_8_reset;
  wire  RetimeWrapper_8_io_flow;
  wire  RetimeWrapper_8_io_in;
  wire  RetimeWrapper_8_io_out;
  wire  _T_2300;
  wire  _T_2302;
  wire  _T_2303;
  wire  RetimeWrapper_9_clock;
  wire  RetimeWrapper_9_reset;
  wire  RetimeWrapper_9_io_flow;
  wire  RetimeWrapper_9_io_in;
  wire  RetimeWrapper_9_io_out;
  wire  _T_2307;
  wire  _T_2309;
  wire  _T_2310;
  wire  RetimeWrapper_10_clock;
  wire  RetimeWrapper_10_reset;
  wire  RetimeWrapper_10_io_flow;
  wire  RetimeWrapper_10_io_in;
  wire  RetimeWrapper_10_io_out;
  wire  _T_2314;
  wire  _T_2316;
  wire  RetimeWrapper_11_clock;
  wire  RetimeWrapper_11_reset;
  wire  RetimeWrapper_11_io_flow;
  wire  RetimeWrapper_11_io_in;
  wire  RetimeWrapper_11_io_out;
  wire  _T_2320;
  wire  _T_2322;
  wire  _T_2323;
  wire  RetimeWrapper_12_clock;
  wire  RetimeWrapper_12_reset;
  wire  RetimeWrapper_12_io_flow;
  wire  RetimeWrapper_12_io_in;
  wire  RetimeWrapper_12_io_out;
  wire  _T_2327;
  wire  _T_2329;
  wire  _T_2330;
  wire  RetimeWrapper_13_clock;
  wire  RetimeWrapper_13_reset;
  wire  RetimeWrapper_13_io_flow;
  wire  RetimeWrapper_13_io_in;
  wire  RetimeWrapper_13_io_out;
  wire  _T_2334;
  wire  _T_2336;
  wire  RetimeWrapper_14_clock;
  wire  RetimeWrapper_14_reset;
  wire  RetimeWrapper_14_io_flow;
  wire  RetimeWrapper_14_io_in;
  wire  RetimeWrapper_14_io_out;
  wire  _T_2340;
  wire  _T_2342;
  wire  _T_2343;
  wire  RetimeWrapper_15_clock;
  wire  RetimeWrapper_15_reset;
  wire  RetimeWrapper_15_io_flow;
  wire  RetimeWrapper_15_io_in;
  wire  RetimeWrapper_15_io_out;
  wire  _T_2347;
  wire  _T_2349;
  wire  _T_2350;
  wire  RetimeWrapper_16_clock;
  wire  RetimeWrapper_16_reset;
  wire  RetimeWrapper_16_io_flow;
  wire  RetimeWrapper_16_io_in;
  wire  RetimeWrapper_16_io_out;
  wire  _T_2354;
  wire  _T_2356;
  wire  RetimeWrapper_17_clock;
  wire  RetimeWrapper_17_reset;
  wire  RetimeWrapper_17_io_flow;
  wire  RetimeWrapper_17_io_in;
  wire  RetimeWrapper_17_io_out;
  wire  _T_2360;
  wire  _T_2362;
  wire  _T_2363;
  wire  RetimeWrapper_18_clock;
  wire  RetimeWrapper_18_reset;
  wire  RetimeWrapper_18_io_flow;
  wire  RetimeWrapper_18_io_in;
  wire  RetimeWrapper_18_io_out;
  wire  _T_2367;
  wire  _T_2369;
  wire  _T_2370;
  wire  RetimeWrapper_19_clock;
  wire  RetimeWrapper_19_reset;
  wire  RetimeWrapper_19_io_flow;
  wire  RetimeWrapper_19_io_in;
  wire  RetimeWrapper_19_io_out;
  wire  _T_2374;
  wire  _T_2376;
  wire  RetimeWrapper_20_clock;
  wire  RetimeWrapper_20_reset;
  wire  RetimeWrapper_20_io_flow;
  wire  RetimeWrapper_20_io_in;
  wire  RetimeWrapper_20_io_out;
  wire  _T_2380;
  wire  RetimeWrapper_21_clock;
  wire  RetimeWrapper_21_reset;
  wire  RetimeWrapper_21_io_flow;
  wire  RetimeWrapper_21_io_in;
  wire  RetimeWrapper_21_io_out;
  wire  _T_2387;
  wire  RetimeWrapper_22_clock;
  wire  RetimeWrapper_22_reset;
  wire  RetimeWrapper_22_io_flow;
  wire  RetimeWrapper_22_io_in;
  wire  RetimeWrapper_22_io_out;
  wire  _T_2394;
  wire  _T_2396;
  wire [31:0] _T_2398_number;
  wire [31:0] _T_2408;
  wire  _T_2423;
  wire  _T_2424;
  wire  _T_2426;
  wire  _T_2429;
  wire  _T_2430;
  reg  _T_2433;
  reg [31:0] _RAND_2;
  wire  _T_2439;
  wire  _T_2441;
  wire  _T_2442;
  wire  _T_2443;
  wire  _T_2444;
  wire  _T_2445;
  reg  _T_2448;
  reg [31:0] _RAND_3;
  wire  _T_2454;
  wire  RetimeWrapper_23_clock;
  wire  RetimeWrapper_23_reset;
  wire  RetimeWrapper_23_io_flow;
  wire  RetimeWrapper_23_io_in;
  wire  RetimeWrapper_23_io_out;
  wire  _T_2458;
  wire  _T_2460;
  wire  RetimeWrapper_24_clock;
  wire  RetimeWrapper_24_reset;
  wire  RetimeWrapper_24_io_flow;
  wire  RetimeWrapper_24_io_in;
  wire  RetimeWrapper_24_io_out;
  wire  _T_2466;
  wire  _T_2468;
  wire  RetimeWrapper_25_clock;
  wire  RetimeWrapper_25_reset;
  wire  RetimeWrapper_25_io_flow;
  wire  RetimeWrapper_25_io_in;
  wire  RetimeWrapper_25_io_out;
  wire  _T_2476;
  wire  _T_2478;
  wire  RetimeWrapper_26_clock;
  wire  RetimeWrapper_26_reset;
  wire  RetimeWrapper_26_io_flow;
  wire  RetimeWrapper_26_io_in;
  wire  RetimeWrapper_26_io_out;
  wire  _T_2483;
  wire  _T_2485;
  wire  _T_2486;
  wire  RetimeWrapper_27_clock;
  wire  RetimeWrapper_27_reset;
  wire  RetimeWrapper_27_io_flow;
  wire  RetimeWrapper_27_io_in;
  wire  RetimeWrapper_27_io_out;
  wire  _T_2490;
  wire  _T_2492;
  wire  RetimeWrapper_28_clock;
  wire  RetimeWrapper_28_reset;
  wire  RetimeWrapper_28_io_flow;
  wire  RetimeWrapper_28_io_in;
  wire  RetimeWrapper_28_io_out;
  wire  _T_2496;
  wire  _T_2498;
  wire  RetimeWrapper_29_clock;
  wire  RetimeWrapper_29_reset;
  wire  RetimeWrapper_29_io_flow;
  wire  RetimeWrapper_29_io_in;
  wire  RetimeWrapper_29_io_out;
  wire  _T_2503;
  wire  _T_2505;
  wire  _T_2506;
  wire  RetimeWrapper_30_clock;
  wire  RetimeWrapper_30_reset;
  wire  RetimeWrapper_30_io_flow;
  wire  RetimeWrapper_30_io_in;
  wire  RetimeWrapper_30_io_out;
  wire  _T_2510;
  wire  _T_2512;
  wire  done_latch_clock;
  wire  done_latch_reset;
  wire  done_latch_io_input_set;
  wire  done_latch_io_input_reset;
  wire  done_latch_io_input_asyn_reset;
  wire  done_latch_io_output_data;
  wire [31:0] _T_2513;
  wire [31:0] _T_2514;
  wire  _T_2517;
  wire  _T_2520;
  wire  _T_2521;
  reg  _T_2524;
  reg [31:0] _RAND_4;
  wire  _T_2530;
  wire  RetimeWrapper_31_clock;
  wire  RetimeWrapper_31_reset;
  wire  RetimeWrapper_31_io_flow;
  wire  RetimeWrapper_31_io_in;
  wire  RetimeWrapper_31_io_out;
  wire  _T_2541;
  wire  _T_2543;
  wire  RetimeWrapper_32_clock;
  wire  RetimeWrapper_32_reset;
  wire  RetimeWrapper_32_io_flow;
  wire  RetimeWrapper_32_io_in;
  wire  RetimeWrapper_32_io_out;
  wire  _T_2549;
  wire  _T_2551;
  wire  _T_2552;
  wire  RetimeWrapper_33_clock;
  wire  RetimeWrapper_33_reset;
  wire  RetimeWrapper_33_io_flow;
  wire  RetimeWrapper_33_io_in;
  wire  RetimeWrapper_33_io_out;
  wire  _T_2556;
  wire  _T_2558;
  wire  _T_2559;
  wire  RetimeWrapper_34_clock;
  wire  RetimeWrapper_34_reset;
  wire  RetimeWrapper_34_io_flow;
  wire  RetimeWrapper_34_io_in;
  wire  RetimeWrapper_34_io_out;
  wire  _T_2563;
  wire  _T_2565;
  wire  RetimeWrapper_35_clock;
  wire  RetimeWrapper_35_reset;
  wire  RetimeWrapper_35_io_flow;
  wire  RetimeWrapper_35_io_in;
  wire  RetimeWrapper_35_io_out;
  wire  _T_2569;
  wire  _T_2571;
  wire  _T_2572;
  wire  RetimeWrapper_36_clock;
  wire  RetimeWrapper_36_reset;
  wire  RetimeWrapper_36_io_flow;
  wire  RetimeWrapper_36_io_in;
  wire  RetimeWrapper_36_io_out;
  wire  _T_2576;
  wire  _T_2578;
  wire  _T_2579;
  wire  RetimeWrapper_37_clock;
  wire  RetimeWrapper_37_reset;
  wire  RetimeWrapper_37_io_flow;
  wire  RetimeWrapper_37_io_in;
  wire  RetimeWrapper_37_io_out;
  wire  _T_2583;
  wire  _T_2585;
  wire  _T_2587;
  wire  _T_2590;
  wire  _T_2591;
  reg  _T_2594;
  reg [31:0] _RAND_5;
  wire  _T_2600;
  wire  RetimeWrapper_38_clock;
  wire  RetimeWrapper_38_reset;
  wire  RetimeWrapper_38_io_flow;
  wire  RetimeWrapper_38_io_in;
  wire  RetimeWrapper_38_io_out;
  wire  _T_2611;
  wire  _T_2613;
  wire  RetimeWrapper_39_clock;
  wire  RetimeWrapper_39_reset;
  wire  RetimeWrapper_39_io_flow;
  wire  RetimeWrapper_39_io_in;
  wire  RetimeWrapper_39_io_out;
  wire  _T_2619;
  wire  _T_2621;
  wire  _T_2622;
  wire  RetimeWrapper_40_clock;
  wire  RetimeWrapper_40_reset;
  wire  RetimeWrapper_40_io_flow;
  wire  RetimeWrapper_40_io_in;
  wire  RetimeWrapper_40_io_out;
  wire  _T_2626;
  wire  _T_2628;
  wire  _T_2629;
  wire  RetimeWrapper_41_clock;
  wire  RetimeWrapper_41_reset;
  wire  RetimeWrapper_41_io_flow;
  wire  RetimeWrapper_41_io_in;
  wire  RetimeWrapper_41_io_out;
  wire  _T_2633;
  wire  _T_2635;
  wire  RetimeWrapper_42_clock;
  wire  RetimeWrapper_42_reset;
  wire  RetimeWrapper_42_io_flow;
  wire  RetimeWrapper_42_io_in;
  wire  RetimeWrapper_42_io_out;
  wire  _T_2639;
  wire  _T_2641;
  wire  _T_2642;
  wire  RetimeWrapper_43_clock;
  wire  RetimeWrapper_43_reset;
  wire  RetimeWrapper_43_io_flow;
  wire  RetimeWrapper_43_io_in;
  wire  RetimeWrapper_43_io_out;
  wire  _T_2646;
  wire  _T_2648;
  wire  _T_2649;
  wire  RetimeWrapper_44_clock;
  wire  RetimeWrapper_44_reset;
  wire  RetimeWrapper_44_io_flow;
  wire  RetimeWrapper_44_io_in;
  wire  RetimeWrapper_44_io_out;
  wire  _T_2653;
  wire  _T_2655;
  wire  _T_2657;
  wire  _T_2660;
  wire  _T_2661;
  reg  _T_2664;
  reg [31:0] _RAND_6;
  wire  _T_2670;
  wire  RetimeWrapper_45_clock;
  wire  RetimeWrapper_45_reset;
  wire  RetimeWrapper_45_io_flow;
  wire  RetimeWrapper_45_io_in;
  wire  RetimeWrapper_45_io_out;
  wire  _T_2681;
  wire  _T_2683;
  wire  RetimeWrapper_46_clock;
  wire  RetimeWrapper_46_reset;
  wire  RetimeWrapper_46_io_flow;
  wire  RetimeWrapper_46_io_in;
  wire  RetimeWrapper_46_io_out;
  wire  _T_2689;
  wire  _T_2691;
  wire  _T_2692;
  wire  RetimeWrapper_47_clock;
  wire  RetimeWrapper_47_reset;
  wire  RetimeWrapper_47_io_flow;
  wire  RetimeWrapper_47_io_in;
  wire  RetimeWrapper_47_io_out;
  wire  _T_2696;
  wire  _T_2698;
  wire  _T_2699;
  wire  RetimeWrapper_48_clock;
  wire  RetimeWrapper_48_reset;
  wire  RetimeWrapper_48_io_flow;
  wire  RetimeWrapper_48_io_in;
  wire  RetimeWrapper_48_io_out;
  wire  _T_2703;
  wire  _T_2705;
  wire  RetimeWrapper_49_clock;
  wire  RetimeWrapper_49_reset;
  wire  RetimeWrapper_49_io_flow;
  wire  RetimeWrapper_49_io_in;
  wire  RetimeWrapper_49_io_out;
  wire  _T_2709;
  wire  _T_2711;
  wire  _T_2712;
  wire  RetimeWrapper_50_clock;
  wire  RetimeWrapper_50_reset;
  wire  RetimeWrapper_50_io_flow;
  wire  RetimeWrapper_50_io_in;
  wire  RetimeWrapper_50_io_out;
  wire  _T_2716;
  wire  _T_2718;
  wire  _T_2719;
  wire  RetimeWrapper_51_clock;
  wire  RetimeWrapper_51_reset;
  wire  RetimeWrapper_51_io_flow;
  wire  RetimeWrapper_51_io_in;
  wire  RetimeWrapper_51_io_out;
  wire  _T_2723;
  wire  _T_2725;
  wire  _T_2729;
  wire  _T_2732;
  wire  _T_2733;
  reg  _T_2736;
  reg [31:0] _RAND_7;
  wire  _T_2742;
  wire  RetimeWrapper_52_clock;
  wire  RetimeWrapper_52_reset;
  wire  RetimeWrapper_52_io_flow;
  wire  RetimeWrapper_52_io_in;
  wire  RetimeWrapper_52_io_out;
  wire  _T_2753;
  wire  _T_2755;
  wire  RetimeWrapper_53_clock;
  wire  RetimeWrapper_53_reset;
  wire  RetimeWrapper_53_io_flow;
  wire  RetimeWrapper_53_io_in;
  wire  RetimeWrapper_53_io_out;
  wire  _T_2761;
  wire  _T_2763;
  wire  _T_2764;
  wire  RetimeWrapper_54_clock;
  wire  RetimeWrapper_54_reset;
  wire  RetimeWrapper_54_io_flow;
  wire  RetimeWrapper_54_io_in;
  wire  RetimeWrapper_54_io_out;
  wire  _T_2768;
  wire  _T_2770;
  wire  _T_2771;
  wire  RetimeWrapper_55_clock;
  wire  RetimeWrapper_55_reset;
  wire  RetimeWrapper_55_io_flow;
  wire  RetimeWrapper_55_io_in;
  wire  RetimeWrapper_55_io_out;
  wire  _T_2775;
  wire  _T_2777;
  wire  RetimeWrapper_56_clock;
  wire  RetimeWrapper_56_reset;
  wire  RetimeWrapper_56_io_flow;
  wire  RetimeWrapper_56_io_in;
  wire  RetimeWrapper_56_io_out;
  wire  _T_2781;
  wire  _T_2783;
  wire  _T_2784;
  wire  RetimeWrapper_57_clock;
  wire  RetimeWrapper_57_reset;
  wire  RetimeWrapper_57_io_flow;
  wire  RetimeWrapper_57_io_in;
  wire  RetimeWrapper_57_io_out;
  wire  _T_2788;
  wire  _T_2790;
  wire  _T_2791;
  wire  RetimeWrapper_58_clock;
  wire  RetimeWrapper_58_reset;
  wire  RetimeWrapper_58_io_flow;
  wire  RetimeWrapper_58_io_in;
  wire  RetimeWrapper_58_io_out;
  wire  _T_2795;
  wire  _T_2797;
  wire  _T_2799;
  wire  _T_2802;
  wire  _T_2803;
  reg  _T_2806;
  reg [31:0] _RAND_8;
  wire  _T_2812;
  wire  _T_2818;
  reg  _T_2821;
  reg [31:0] _RAND_9;
  wire  _T_2827;
  wire  RetimeWrapper_59_clock;
  wire  RetimeWrapper_59_reset;
  wire  RetimeWrapper_59_io_flow;
  wire  RetimeWrapper_59_io_in;
  wire  RetimeWrapper_59_io_out;
  wire  _T_2831;
  wire  _T_2833;
  wire  RetimeWrapper_60_clock;
  wire  RetimeWrapper_60_reset;
  wire  RetimeWrapper_60_io_flow;
  wire  RetimeWrapper_60_io_in;
  wire  RetimeWrapper_60_io_out;
  wire  _T_2846;
  wire  _T_2848;
  wire  RetimeWrapper_61_clock;
  wire  RetimeWrapper_61_reset;
  wire  RetimeWrapper_61_io_flow;
  wire  RetimeWrapper_61_io_in;
  wire  RetimeWrapper_61_io_out;
  wire  _T_2859;
  wire  _T_2861;
  wire  RetimeWrapper_62_clock;
  wire  RetimeWrapper_62_reset;
  wire  RetimeWrapper_62_io_flow;
  wire  RetimeWrapper_62_io_in;
  wire  RetimeWrapper_62_io_out;
  wire  _T_2867;
  wire  _T_2869;
  wire  _T_2870;
  wire  RetimeWrapper_63_clock;
  wire  RetimeWrapper_63_reset;
  wire  RetimeWrapper_63_io_flow;
  wire  RetimeWrapper_63_io_in;
  wire  RetimeWrapper_63_io_out;
  wire  _T_2874;
  wire  _T_2876;
  wire  _T_2877;
  wire  _T_2878;
  wire  _T_2879;
  wire  RetimeWrapper_64_clock;
  wire  RetimeWrapper_64_reset;
  wire  RetimeWrapper_64_io_flow;
  wire  RetimeWrapper_64_io_in;
  wire  RetimeWrapper_64_io_out;
  wire  _T_2883;
  wire  _T_2885;
  wire  _T_2886;
  wire  _T_2887;
  wire  _T_2888;
  wire  RetimeWrapper_65_clock;
  wire  RetimeWrapper_65_reset;
  wire  RetimeWrapper_65_io_flow;
  wire  RetimeWrapper_65_io_in;
  wire  RetimeWrapper_65_io_out;
  wire  _T_2892;
  wire  _T_2894;
  wire  RetimeWrapper_66_clock;
  wire  RetimeWrapper_66_reset;
  wire  RetimeWrapper_66_io_flow;
  wire  RetimeWrapper_66_io_in;
  wire  RetimeWrapper_66_io_out;
  wire  _T_2898;
  wire  _T_2900;
  wire  _T_2901;
  wire  RetimeWrapper_67_clock;
  wire  RetimeWrapper_67_reset;
  wire  RetimeWrapper_67_io_flow;
  wire  RetimeWrapper_67_io_in;
  wire  RetimeWrapper_67_io_out;
  wire  _T_2905;
  wire  _T_2907;
  wire  _T_2908;
  wire  RetimeWrapper_68_clock;
  wire  RetimeWrapper_68_reset;
  wire  RetimeWrapper_68_io_flow;
  wire  RetimeWrapper_68_io_in;
  wire  RetimeWrapper_68_io_out;
  wire  _T_2912;
  wire  _T_2914;
  wire  _T_2915;
  wire  _T_2917;
  wire  RetimeWrapper_69_clock;
  wire  RetimeWrapper_69_reset;
  wire  RetimeWrapper_69_io_flow;
  wire  RetimeWrapper_69_io_in;
  wire  RetimeWrapper_69_io_out;
  wire  _T_2928;
  wire  _T_2930;
  wire  RetimeWrapper_70_clock;
  wire  RetimeWrapper_70_reset;
  wire  RetimeWrapper_70_io_flow;
  wire  RetimeWrapper_70_io_in;
  wire  RetimeWrapper_70_io_out;
  wire  _T_2936;
  wire  _T_2938;
  wire  _T_2939;
  wire  RetimeWrapper_71_clock;
  wire  RetimeWrapper_71_reset;
  wire  RetimeWrapper_71_io_flow;
  wire  RetimeWrapper_71_io_in;
  wire  RetimeWrapper_71_io_out;
  wire  _T_2943;
  wire  _T_2945;
  wire  _T_2946;
  wire  _T_2947;
  wire  _T_2948;
  wire  RetimeWrapper_72_clock;
  wire  RetimeWrapper_72_reset;
  wire  RetimeWrapper_72_io_flow;
  wire  RetimeWrapper_72_io_in;
  wire  RetimeWrapper_72_io_out;
  wire  _T_2952;
  wire  _T_2954;
  wire  _T_2955;
  wire  _T_2956;
  wire  _T_2957;
  wire  RetimeWrapper_73_clock;
  wire  RetimeWrapper_73_reset;
  wire  RetimeWrapper_73_io_flow;
  wire  RetimeWrapper_73_io_in;
  wire  RetimeWrapper_73_io_out;
  wire  _T_2961;
  wire  _T_2963;
  wire  RetimeWrapper_74_clock;
  wire  RetimeWrapper_74_reset;
  wire  RetimeWrapper_74_io_flow;
  wire  RetimeWrapper_74_io_in;
  wire  RetimeWrapper_74_io_out;
  wire  _T_2967;
  wire  _T_2969;
  wire  _T_2970;
  wire  RetimeWrapper_75_clock;
  wire  RetimeWrapper_75_reset;
  wire  RetimeWrapper_75_io_flow;
  wire  RetimeWrapper_75_io_in;
  wire  RetimeWrapper_75_io_out;
  wire  _T_2974;
  wire  _T_2976;
  wire  _T_2977;
  wire  RetimeWrapper_76_clock;
  wire  RetimeWrapper_76_reset;
  wire  RetimeWrapper_76_io_flow;
  wire  RetimeWrapper_76_io_in;
  wire  RetimeWrapper_76_io_out;
  wire  _T_2981;
  wire  _T_2983;
  wire  _T_2984;
  wire  _T_2986;
  wire  _T_2987;
  wire  _T_2990;
  wire  _T_2991;
  wire  _T_2992;
  wire  _T_2993;
  reg  _T_2996;
  reg [31:0] _RAND_10;
  wire  _T_3002;
  wire  RetimeWrapper_77_clock;
  wire  RetimeWrapper_77_reset;
  wire  RetimeWrapper_77_io_flow;
  wire  RetimeWrapper_77_io_in;
  wire  RetimeWrapper_77_io_out;
  wire  _T_3007;
  wire  _T_3009;
  wire  RetimeWrapper_78_clock;
  wire  RetimeWrapper_78_reset;
  wire  RetimeWrapper_78_io_flow;
  wire  RetimeWrapper_78_io_in;
  wire  RetimeWrapper_78_io_out;
  wire  _T_3016;
  wire  _T_3018;
  wire  _T_3025;
  wire [63:0] _T_3026;
  wire [31:0] _T_3027;
  wire  _T_3028;
  wire  _T_3029;
  wire  _T_3034;
  wire  _T_3035;
  wire  _T_3037;
  wire  RetimeWrapper_79_clock;
  wire  RetimeWrapper_79_reset;
  wire  RetimeWrapper_79_io_flow;
  wire  RetimeWrapper_79_io_in;
  wire  RetimeWrapper_79_io_out;
  wire  _T_3048;
  wire  _T_3050;
  wire  RetimeWrapper_80_clock;
  wire  RetimeWrapper_80_reset;
  wire  RetimeWrapper_80_io_flow;
  wire  RetimeWrapper_80_io_in;
  wire  RetimeWrapper_80_io_out;
  wire  _T_3056;
  wire  _T_3058;
  wire  _T_3059;
  wire  RetimeWrapper_81_clock;
  wire  RetimeWrapper_81_reset;
  wire  RetimeWrapper_81_io_flow;
  wire  RetimeWrapper_81_io_in;
  wire  RetimeWrapper_81_io_out;
  wire  _T_3063;
  wire  _T_3065;
  wire  _T_3066;
  wire  _T_3067;
  wire  RetimeWrapper_82_clock;
  wire  RetimeWrapper_82_reset;
  wire  RetimeWrapper_82_io_flow;
  wire  RetimeWrapper_82_io_in;
  wire  RetimeWrapper_82_io_out;
  wire  _T_3071;
  wire  _T_3073;
  wire  _T_3075;
  wire  _T_3076;
  wire  RetimeWrapper_83_clock;
  wire  RetimeWrapper_83_reset;
  wire  RetimeWrapper_83_io_flow;
  wire  RetimeWrapper_83_io_in;
  wire  RetimeWrapper_83_io_out;
  wire  _T_3080;
  wire  _T_3082;
  wire  RetimeWrapper_84_clock;
  wire  RetimeWrapper_84_reset;
  wire  RetimeWrapper_84_io_flow;
  wire  RetimeWrapper_84_io_in;
  wire  RetimeWrapper_84_io_out;
  wire  _T_3086;
  wire  _T_3088;
  wire  _T_3089;
  wire  RetimeWrapper_85_clock;
  wire  RetimeWrapper_85_reset;
  wire  RetimeWrapper_85_io_flow;
  wire  RetimeWrapper_85_io_in;
  wire  RetimeWrapper_85_io_out;
  wire  _T_3093;
  wire  _T_3095;
  wire  _T_3096;
  wire  _T_3097;
  wire  RetimeWrapper_86_clock;
  wire  RetimeWrapper_86_reset;
  wire  RetimeWrapper_86_io_flow;
  wire  RetimeWrapper_86_io_in;
  wire  RetimeWrapper_86_io_out;
  wire  _T_3104;
  wire  _T_3106;
  wire  _T_3109;
  wire  _T_3110;
  wire  _T_3111;
  wire  _T_3112;
  reg  _T_3115;
  reg [31:0] _RAND_11;
  wire  _T_3121;
  wire  RetimeWrapper_87_clock;
  wire  RetimeWrapper_87_reset;
  wire  RetimeWrapper_87_io_flow;
  wire  RetimeWrapper_87_io_in;
  wire  RetimeWrapper_87_io_out;
  wire  _T_3125;
  wire  _T_3127;
  wire  RetimeWrapper_88_clock;
  wire  RetimeWrapper_88_reset;
  wire  RetimeWrapper_88_io_flow;
  wire  RetimeWrapper_88_io_in;
  wire  RetimeWrapper_88_io_out;
  wire  _T_3133;
  wire  _T_3135;
  wire [31:0] _T_3139;
  wire  _T_3408;
  wire  _T_3410;
  wire  _T_3411;
  wire  _T_3412;
  wire  RetimeWrapper_89_clock;
  wire  RetimeWrapper_89_reset;
  wire  RetimeWrapper_89_io_flow;
  wire  RetimeWrapper_89_io_in;
  wire  RetimeWrapper_89_io_out;
  wire  _T_3419;
  wire  _T_3421;
  wire  RetimeWrapper_90_clock;
  wire  RetimeWrapper_90_reset;
  wire  RetimeWrapper_90_io_flow;
  wire  RetimeWrapper_90_io_in;
  wire  RetimeWrapper_90_io_out;
  wire  _T_3425;
  wire  _T_3427;
  wire [31:0] _T_3504_number;
  wire [31:0] _T_3506_number;
  wire [31:0] _T_3514;
  wire [31:0] _T_3525;
  wire [31:0] _T_3529;
  wire [31:0] _T_3530;
  wire  _T_3531;
  wire  RetimeWrapper_91_clock;
  wire  RetimeWrapper_91_reset;
  wire  RetimeWrapper_91_io_flow;
  wire  RetimeWrapper_91_io_in;
  wire  RetimeWrapper_91_io_out;
  wire  _T_3565;
  wire  _T_3567;
  wire [31:0] _T_3569_number;
  wire [31:0] _T_3579;
  wire  _T_3594;
  wire  _T_3595;
  wire  _T_3596;
  wire  _T_3598;
  wire  RetimeWrapper_92_clock;
  wire  RetimeWrapper_92_reset;
  wire  RetimeWrapper_92_io_flow;
  wire  RetimeWrapper_92_io_in;
  wire  RetimeWrapper_92_io_out;
  wire  _T_3609;
  wire  _T_3611;
  wire  RetimeWrapper_93_clock;
  wire  RetimeWrapper_93_reset;
  wire  RetimeWrapper_93_io_flow;
  wire  RetimeWrapper_93_io_in;
  wire  RetimeWrapper_93_io_out;
  wire  _T_3617;
  wire  _T_3619;
  wire  _T_3620;
  wire  RetimeWrapper_94_clock;
  wire  RetimeWrapper_94_reset;
  wire  RetimeWrapper_94_io_flow;
  wire  RetimeWrapper_94_io_in;
  wire  RetimeWrapper_94_io_out;
  wire  _T_3624;
  wire  _T_3626;
  wire  _T_3627;
  wire  _T_3628;
  wire  _T_3629;
  wire  RetimeWrapper_95_clock;
  wire  RetimeWrapper_95_reset;
  wire  RetimeWrapper_95_io_flow;
  wire  RetimeWrapper_95_io_in;
  wire  RetimeWrapper_95_io_out;
  wire  _T_3633;
  wire  _T_3635;
  wire  _T_3636;
  wire  _T_3637;
  wire  _T_3638;
  wire  RetimeWrapper_96_clock;
  wire  RetimeWrapper_96_reset;
  wire  RetimeWrapper_96_io_flow;
  wire  RetimeWrapper_96_io_in;
  wire  RetimeWrapper_96_io_out;
  wire  _T_3642;
  wire  _T_3644;
  wire  RetimeWrapper_97_clock;
  wire  RetimeWrapper_97_reset;
  wire  RetimeWrapper_97_io_flow;
  wire  RetimeWrapper_97_io_in;
  wire  RetimeWrapper_97_io_out;
  wire  _T_3648;
  wire  _T_3650;
  wire  _T_3651;
  wire  RetimeWrapper_98_clock;
  wire  RetimeWrapper_98_reset;
  wire  RetimeWrapper_98_io_flow;
  wire  RetimeWrapper_98_io_in;
  wire  RetimeWrapper_98_io_out;
  wire  _T_3655;
  wire  _T_3657;
  wire  _T_3658;
  wire  RetimeWrapper_99_clock;
  wire  RetimeWrapper_99_reset;
  wire  RetimeWrapper_99_io_flow;
  wire  RetimeWrapper_99_io_in;
  wire  RetimeWrapper_99_io_out;
  wire  _T_3662;
  wire  _T_3664;
  wire  _T_3665;
  wire  _T_3667;
  wire  RetimeWrapper_100_clock;
  wire  RetimeWrapper_100_reset;
  wire  RetimeWrapper_100_io_flow;
  wire  RetimeWrapper_100_io_in;
  wire  RetimeWrapper_100_io_out;
  wire  _T_3678;
  wire  _T_3680;
  wire  RetimeWrapper_101_clock;
  wire  RetimeWrapper_101_reset;
  wire  RetimeWrapper_101_io_flow;
  wire  RetimeWrapper_101_io_in;
  wire  RetimeWrapper_101_io_out;
  wire  _T_3686;
  wire  _T_3688;
  wire  _T_3689;
  wire  RetimeWrapper_102_clock;
  wire  RetimeWrapper_102_reset;
  wire  RetimeWrapper_102_io_flow;
  wire  RetimeWrapper_102_io_in;
  wire  RetimeWrapper_102_io_out;
  wire  _T_3693;
  wire  _T_3695;
  wire  _T_3696;
  wire  _T_3697;
  wire  _T_3698;
  wire  RetimeWrapper_103_clock;
  wire  RetimeWrapper_103_reset;
  wire  RetimeWrapper_103_io_flow;
  wire  RetimeWrapper_103_io_in;
  wire  RetimeWrapper_103_io_out;
  wire  _T_3702;
  wire  _T_3704;
  wire  _T_3705;
  wire  _T_3706;
  wire  _T_3707;
  wire  RetimeWrapper_104_clock;
  wire  RetimeWrapper_104_reset;
  wire  RetimeWrapper_104_io_flow;
  wire  RetimeWrapper_104_io_in;
  wire  RetimeWrapper_104_io_out;
  wire  _T_3711;
  wire  _T_3713;
  wire  RetimeWrapper_105_clock;
  wire  RetimeWrapper_105_reset;
  wire  RetimeWrapper_105_io_flow;
  wire  RetimeWrapper_105_io_in;
  wire  RetimeWrapper_105_io_out;
  wire  _T_3717;
  wire  _T_3719;
  wire  _T_3720;
  wire  RetimeWrapper_106_clock;
  wire  RetimeWrapper_106_reset;
  wire  RetimeWrapper_106_io_flow;
  wire  RetimeWrapper_106_io_in;
  wire  RetimeWrapper_106_io_out;
  wire  _T_3724;
  wire  _T_3726;
  wire  _T_3727;
  wire  RetimeWrapper_107_clock;
  wire  RetimeWrapper_107_reset;
  wire  RetimeWrapper_107_io_flow;
  wire  RetimeWrapper_107_io_in;
  wire  RetimeWrapper_107_io_out;
  wire  _T_3731;
  wire  _T_3733;
  wire  _T_3734;
  wire  _T_3736;
  wire  _T_3737;
  wire  _T_3740;
  wire  _T_3741;
  wire  _T_3742;
  wire  _T_3743;
  reg  _T_3746;
  reg [31:0] _RAND_12;
  wire  _T_3752;
  wire  RetimeWrapper_108_clock;
  wire  RetimeWrapper_108_reset;
  wire  RetimeWrapper_108_io_flow;
  wire  RetimeWrapper_108_io_in;
  wire  RetimeWrapper_108_io_out;
  wire  _T_3757;
  wire  _T_3759;
  wire  RetimeWrapper_109_clock;
  wire  RetimeWrapper_109_reset;
  wire  RetimeWrapper_109_io_flow;
  wire  RetimeWrapper_109_io_in;
  wire  RetimeWrapper_109_io_out;
  wire  _T_3766;
  wire  _T_3768;
  wire  _T_3775;
  wire [63:0] _T_3776;
  wire [31:0] _T_3777;
  wire  _T_3778;
  wire  _T_3779;
  wire  _T_3784;
  wire  _T_3785;
  wire  _T_3787;
  wire  RetimeWrapper_110_clock;
  wire  RetimeWrapper_110_reset;
  wire  RetimeWrapper_110_io_flow;
  wire  RetimeWrapper_110_io_in;
  wire  RetimeWrapper_110_io_out;
  wire  _T_3798;
  wire  _T_3800;
  wire  RetimeWrapper_111_clock;
  wire  RetimeWrapper_111_reset;
  wire  RetimeWrapper_111_io_flow;
  wire  RetimeWrapper_111_io_in;
  wire  RetimeWrapper_111_io_out;
  wire  _T_3806;
  wire  _T_3808;
  wire  _T_3809;
  wire  RetimeWrapper_112_clock;
  wire  RetimeWrapper_112_reset;
  wire  RetimeWrapper_112_io_flow;
  wire  RetimeWrapper_112_io_in;
  wire  RetimeWrapper_112_io_out;
  wire  _T_3813;
  wire  _T_3815;
  wire  _T_3816;
  wire  _T_3817;
  wire  RetimeWrapper_113_clock;
  wire  RetimeWrapper_113_reset;
  wire  RetimeWrapper_113_io_flow;
  wire  RetimeWrapper_113_io_in;
  wire  RetimeWrapper_113_io_out;
  wire  _T_3821;
  wire  _T_3823;
  wire  _T_3825;
  wire  _T_3826;
  wire  RetimeWrapper_114_clock;
  wire  RetimeWrapper_114_reset;
  wire  RetimeWrapper_114_io_flow;
  wire  RetimeWrapper_114_io_in;
  wire  RetimeWrapper_114_io_out;
  wire  _T_3830;
  wire  _T_3832;
  wire  RetimeWrapper_115_clock;
  wire  RetimeWrapper_115_reset;
  wire  RetimeWrapper_115_io_flow;
  wire  RetimeWrapper_115_io_in;
  wire  RetimeWrapper_115_io_out;
  wire  _T_3836;
  wire  _T_3838;
  wire  _T_3839;
  wire  RetimeWrapper_116_clock;
  wire  RetimeWrapper_116_reset;
  wire  RetimeWrapper_116_io_flow;
  wire  RetimeWrapper_116_io_in;
  wire  RetimeWrapper_116_io_out;
  wire  _T_3843;
  wire  _T_3845;
  wire  _T_3846;
  wire  _T_3847;
  wire  RetimeWrapper_117_clock;
  wire  RetimeWrapper_117_reset;
  wire  RetimeWrapper_117_io_flow;
  wire  RetimeWrapper_117_io_in;
  wire  RetimeWrapper_117_io_out;
  wire [31:0] _T_3855_number;
  wire [31:0] _T_3857_number;
  wire [31:0] _T_3865;
  wire [31:0] _T_3870_number;
  wire [33:0] _GEN_0;
  wire [33:0] _T_3871;
  wire [5:0] x3181;
  wire [31:0] _T_3873_number;
  wire [33:0] _GEN_1;
  wire [33:0] _T_3874;
  wire [32:0] _T_3876_number;
  wire [32:0] _T_3878_number;
  wire [32:0] _T_3880_number;
  wire [32:0] _T_3888;
  wire  _T_3891;
  wire [32:0] _T_3893;
  wire [32:0] _T_3901;
  wire  _T_3904;
  wire [32:0] _T_3906;
  wire [33:0] _T_3907;
  wire [33:0] _T_3908;
  wire [32:0] _T_3909;
  wire [31:0] _T_3911_number;
  wire [31:0] _T_3925;
  wire [31:0] _T_3929;
  wire [32:0] _T_3931_number;
  wire [32:0] _T_3933_number;
  wire [32:0] _T_3935_number;
  wire [32:0] _T_3943;
  wire [32:0] _T_3956;
  wire  _T_3959;
  wire [32:0] _T_3961;
  wire [33:0] _T_3962;
  wire [32:0] _T_3963;
  wire [31:0] _T_3965_number;
  wire [31:0] _T_3979;
  wire [31:0] _T_3983;
  wire [5:0] x3188;
  wire [31:0] _T_3989_number;
  wire [31:0] _T_3999;
  wire  _T_4014;
  wire [32:0] _T_4020_number;
  wire [32:0] _T_4024_number;
  wire [32:0] _T_4045;
  wire  _T_4048;
  wire [32:0] _T_4050;
  wire [33:0] _T_4051;
  wire [33:0] _T_4052;
  wire [32:0] _T_4053;
  wire [31:0] _T_4055_number;
  wire [31:0] _T_4069;
  wire [31:0] _T_4073;
  wire [31:0] _T_4078;
  wire [31:0] _T_4080_number;
  wire [1:0] _T_4085;
  wire [29:0] _T_4086;
  wire [31:0] _T_4087;
  wire [31:0] _T_4089_number;
  wire  _T_4090;
  wire [1:0] _T_4094;
  wire [29:0] _T_4095;
  wire [31:0] _T_4096;
  wire [32:0] _T_4098_number;
  wire [32:0] _T_4100_number;
  wire [32:0] _T_4102_number;
  wire [32:0] _T_4110;
  wire  _T_4113;
  wire [32:0] _T_4115;
  wire [32:0] _T_4123;
  wire  _T_4126;
  wire [32:0] _T_4128;
  wire [33:0] _T_4129;
  wire [32:0] _T_4130;
  wire [31:0] _T_4132_number;
  wire [31:0] _T_4146;
  wire [31:0] _T_4150;
  wire [32:0] _T_4152_number;
  wire [32:0] _T_4154_number;
  wire [32:0] _T_4156_number;
  wire [32:0] _T_4164;
  wire [32:0] _T_4177;
  wire [33:0] _T_4183;
  wire [32:0] _T_4184;
  wire [31:0] _T_4186_number;
  wire [31:0] _T_4200;
  wire [31:0] _T_4204;
  wire [32:0] _T_4206_number;
  wire [32:0] _T_4208_number;
  wire [32:0] _T_4210_number;
  wire [32:0] _T_4218;
  wire  _T_4221;
  wire [32:0] _T_4223;
  wire [32:0] _T_4231;
  wire  _T_4234;
  wire [32:0] _T_4236;
  wire [33:0] _T_4237;
  wire [32:0] _T_4238;
  wire [31:0] _T_4240_number;
  wire [31:0] _T_4254;
  wire [31:0] _T_4258;
  wire [32:0] _T_4260_number;
  wire [32:0] _T_4262_number;
  wire [32:0] _T_4264_number;
  wire [32:0] _T_4272;
  wire [32:0] _T_4285;
  wire [33:0] _T_4291;
  wire [32:0] _T_4292;
  wire [31:0] _T_4294_number;
  wire [31:0] _T_4308;
  wire [31:0] _T_4312;
  wire [32:0] _T_4314_number;
  wire [32:0] _T_4316_number;
  wire [32:0] _T_4318_number;
  wire [32:0] _T_4326;
  wire  _T_4329;
  wire [32:0] _T_4331;
  wire [32:0] _T_4339;
  wire [32:0] _T_4344;
  wire [33:0] _T_4345;
  wire [32:0] _T_4346;
  wire [31:0] _T_4348_number;
  wire [31:0] _T_4362;
  wire [31:0] _T_4366;
  wire [63:0] _T_4374;
  wire  _T_4377;
  wire [31:0] _T_4381;
  wire [63:0] _T_4383;
  wire [63:0] _T_4385_number;
  wire [63:0] _T_4387_number;
  wire [63:0] _T_4395;
  wire [64:0] _T_4400_number;
  wire [64:0] _T_4402_number;
  wire [64:0] _T_4404_number;
  wire [64:0] _T_4412;
  wire  _T_4415;
  wire [64:0] _T_4417;
  wire [64:0] _T_4425;
  wire  _T_4428;
  wire [64:0] _T_4430;
  wire [65:0] _T_4431;
  wire [64:0] _T_4432;
  wire [63:0] _T_4434_number;
  wire [63:0] _T_4448;
  wire [63:0] _T_4452;
  wire [63:0] _T_4460;
  wire [32:0] _T_4465;
  wire [96:0] _T_4466;
  wire  _T_4472;
  wire  _T_4473;
  wire  _T_4480;
  wire [63:0] _T_4481;
  wire [95:0] _T_4482;
  wire [95:0] _T_4485_0;
  wire  _T_4499_0;
  wire  _T_4503;
  wire  _T_4505;
  wire  _T_4506;
  wire  _T_4509;
  wire  _T_4510;
  wire  _T_4511;
  wire  _T_4512;
  reg  _T_4515;
  reg [31:0] _RAND_13;
  wire  _T_4521;
  wire  RetimeWrapper_118_clock;
  wire  RetimeWrapper_118_reset;
  wire  RetimeWrapper_118_io_flow;
  wire  RetimeWrapper_118_io_in;
  wire  RetimeWrapper_118_io_out;
  wire  _T_4526;
  wire  _T_4528;
  wire  RetimeWrapper_119_clock;
  wire  RetimeWrapper_119_reset;
  wire  RetimeWrapper_119_io_flow;
  wire  RetimeWrapper_119_io_in;
  wire  RetimeWrapper_119_io_out;
  wire  _T_4535;
  wire  _T_4537;
  wire  _T_4544;
  wire [63:0] _T_4545;
  wire [31:0] _T_4546;
  wire  _T_4547;
  wire  _T_4548;
  wire  _T_4553;
  wire  _T_4554;
  wire  _T_4556;
  wire  RetimeWrapper_120_clock;
  wire  RetimeWrapper_120_reset;
  wire  RetimeWrapper_120_io_flow;
  wire  RetimeWrapper_120_io_in;
  wire  RetimeWrapper_120_io_out;
  wire  _T_4567;
  wire  _T_4569;
  wire  RetimeWrapper_121_clock;
  wire  RetimeWrapper_121_reset;
  wire  RetimeWrapper_121_io_flow;
  wire  RetimeWrapper_121_io_in;
  wire  RetimeWrapper_121_io_out;
  wire  _T_4575;
  wire  _T_4577;
  wire  _T_4578;
  wire  RetimeWrapper_122_clock;
  wire  RetimeWrapper_122_reset;
  wire  RetimeWrapper_122_io_flow;
  wire  RetimeWrapper_122_io_in;
  wire  RetimeWrapper_122_io_out;
  wire  _T_4582;
  wire  _T_4584;
  wire  _T_4585;
  wire  _T_4586;
  wire  RetimeWrapper_123_clock;
  wire  RetimeWrapper_123_reset;
  wire  RetimeWrapper_123_io_flow;
  wire  RetimeWrapper_123_io_in;
  wire  RetimeWrapper_123_io_out;
  wire  _T_4590;
  wire  _T_4592;
  wire  _T_4594;
  wire  _T_4595;
  wire  RetimeWrapper_124_clock;
  wire  RetimeWrapper_124_reset;
  wire  RetimeWrapper_124_io_flow;
  wire  RetimeWrapper_124_io_in;
  wire  RetimeWrapper_124_io_out;
  wire  _T_4599;
  wire  _T_4601;
  wire  RetimeWrapper_125_clock;
  wire  RetimeWrapper_125_reset;
  wire  RetimeWrapper_125_io_flow;
  wire  RetimeWrapper_125_io_in;
  wire  RetimeWrapper_125_io_out;
  wire  _T_4605;
  wire  _T_4607;
  wire  _T_4608;
  wire  RetimeWrapper_126_clock;
  wire  RetimeWrapper_126_reset;
  wire  RetimeWrapper_126_io_flow;
  wire  RetimeWrapper_126_io_in;
  wire  RetimeWrapper_126_io_out;
  wire  _T_4612;
  wire  _T_4614;
  wire  _T_4615;
  wire  _T_4616;
  wire  RetimeWrapper_127_clock;
  wire  RetimeWrapper_127_reset;
  wire  RetimeWrapper_127_io_flow;
  wire  RetimeWrapper_127_io_in;
  wire  RetimeWrapper_127_io_out;
  wire  _T_4623;
  wire  _T_4625;
  wire  _T_4628;
  wire  _T_4629;
  wire  _T_4630;
  wire  _T_4631;
  reg  _T_4634;
  reg [31:0] _RAND_14;
  wire  _T_4640;
  wire  RetimeWrapper_128_clock;
  wire  RetimeWrapper_128_reset;
  wire  RetimeWrapper_128_io_flow;
  wire  RetimeWrapper_128_io_in;
  wire  RetimeWrapper_128_io_out;
  wire  _T_4644;
  wire  _T_4646;
  wire  RetimeWrapper_129_clock;
  wire  RetimeWrapper_129_reset;
  wire  RetimeWrapper_129_io_flow;
  wire  RetimeWrapper_129_io_in;
  wire  RetimeWrapper_129_io_out;
  wire  _T_4652;
  wire  _T_4654;
  wire [31:0] _T_4658;
  wire  _T_4927;
  wire  _T_4929;
  wire  _T_4930;
  wire  _T_4931;
  wire  RetimeWrapper_130_clock;
  wire  RetimeWrapper_130_reset;
  wire  RetimeWrapper_130_io_flow;
  wire  RetimeWrapper_130_io_in;
  wire  RetimeWrapper_130_io_out;
  wire  _T_4938;
  wire  _T_4940;
  wire  RetimeWrapper_131_clock;
  wire  RetimeWrapper_131_reset;
  wire  RetimeWrapper_131_io_flow;
  wire  RetimeWrapper_131_io_in;
  wire  RetimeWrapper_131_io_out;
  wire  _T_4944;
  wire  _T_4946;
  wire [31:0] _T_5023_number;
  wire [31:0] _T_5025_number;
  wire [31:0] _T_5033;
  wire [31:0] _T_5044;
  wire [31:0] _T_5048;
  wire [31:0] _T_5049;
  wire  _T_5050;
  wire  RetimeWrapper_132_clock;
  wire  RetimeWrapper_132_reset;
  wire  RetimeWrapper_132_io_flow;
  wire  RetimeWrapper_132_io_in;
  wire  RetimeWrapper_132_io_out;
  wire  _T_5084;
  wire  _T_5086;
  wire [31:0] _T_5088_number;
  wire [31:0] _T_5098;
  wire  _T_5113;
  wire  _T_5114;
  wire [31:0] _T_5115;
  wire  _T_5382;
  wire  _T_5385;
  wire  _T_5386;
  reg  _T_5389;
  reg [31:0] _RAND_15;
  wire  _T_5395;
  wire  _T_5397;
  wire  _T_5398;
  wire  _T_5399;
  wire  _T_5400;
  wire  _T_5403;
  wire  RetimeWrapper_133_clock;
  wire  RetimeWrapper_133_reset;
  wire  RetimeWrapper_133_io_flow;
  wire  RetimeWrapper_133_io_in;
  wire  RetimeWrapper_133_io_out;
  wire  _T_5407;
  wire  _T_5409;
  wire  _T_5416;
  wire [31:0] _T_5491_number;
  wire [31:0] _T_5493_number;
  wire [31:0] _T_5501;
  wire [31:0] _T_5512;
  wire [31:0] _T_5516;
  wire [31:0] _T_5517;
  wire  _T_5518;
  wire [31:0] _T_5621_number;
  wire [31:0] _T_5623_number;
  wire [31:0] _T_5631;
  wire [31:0] _T_5642;
  wire [31:0] _T_5646;
  wire [31:0] _T_5647;
  wire  _T_5648;
  wire [31:0] _T_5751_number;
  wire [31:0] _T_5753_number;
  wire [31:0] _T_5761;
  wire [31:0] _T_5772;
  wire [31:0] _T_5776;
  wire [31:0] _T_5777;
  wire  _T_5778;
  wire [31:0] _T_5881_number;
  wire [31:0] _T_5883_number;
  wire [31:0] _T_5891;
  wire [31:0] _T_5902;
  wire [31:0] _T_5906;
  wire [31:0] _T_5907;
  wire  _T_5908;
  wire  RetimeWrapper_134_clock;
  wire  RetimeWrapper_134_reset;
  wire  RetimeWrapper_134_io_flow;
  wire  RetimeWrapper_134_io_in;
  wire  RetimeWrapper_134_io_out;
  wire  _T_5942;
  wire  _T_5944;
  wire [31:0] _T_5946_number;
  wire [31:0] _T_5956;
  wire  _T_5971;
  wire  _T_5972;
  wire [31:0] _T_5973;
  wire  _T_6240;
  wire  _T_6243;
  wire  _T_6244;
  reg  _T_6247;
  reg [31:0] _RAND_16;
  wire  _T_6253;
  wire  _T_6255;
  wire  _T_6256;
  wire  _T_6257;
  wire  _T_6258;
  wire  _T_6261;
  wire  RetimeWrapper_135_clock;
  wire  RetimeWrapper_135_reset;
  wire  RetimeWrapper_135_io_flow;
  wire  RetimeWrapper_135_io_in;
  wire  RetimeWrapper_135_io_out;
  wire  _T_6265;
  wire  _T_6267;
  wire  _T_6274;
  wire [31:0] _T_6349_number;
  wire [31:0] _T_6351_number;
  wire [31:0] _T_6359;
  wire [31:0] _T_6370;
  wire [31:0] _T_6374;
  wire [31:0] _T_6375;
  wire  _T_6376;
  wire [31:0] _T_6479_number;
  wire [31:0] _T_6481_number;
  wire [31:0] _T_6489;
  wire [31:0] _T_6500;
  wire [31:0] _T_6504;
  wire [31:0] _T_6505;
  wire  _T_6506;
  wire [31:0] _T_6609_number;
  wire [31:0] _T_6611_number;
  wire [31:0] _T_6619;
  wire [31:0] _T_6630;
  wire [31:0] _T_6634;
  wire [31:0] _T_6635;
  wire  _T_6636;
  wire [31:0] _T_6739_number;
  wire [31:0] _T_6741_number;
  wire [31:0] _T_6749;
  wire [31:0] _T_6760;
  wire [31:0] _T_6764;
  wire [31:0] _T_6765;
  wire  _T_6766;
  wire  RetimeWrapper_136_clock;
  wire  RetimeWrapper_136_reset;
  wire  RetimeWrapper_136_io_flow;
  wire  RetimeWrapper_136_io_in;
  wire  RetimeWrapper_136_io_out;
  wire  _T_6800;
  wire  _T_6802;
  wire [31:0] _T_6804_number;
  wire [31:0] _T_6814;
  wire  _T_6829;
  wire  _T_6830;
  wire [32:0] _T_6832_number;
  wire [32:0] _T_6834_number;
  wire [32:0] _T_6836_number;
  wire [7:0] _T_6840;
  wire [7:0] _T_6842;
  wire [24:0] _T_6844;
  wire [7:0] _T_6845;
  wire  _T_6846;
  wire [23:0] _T_6847;
  wire [24:0] _T_6848;
  wire [32:0] _T_6849;
  wire [7:0] _T_6853;
  wire [7:0] _T_6855;
  wire [24:0] _T_6857;
  wire [7:0] _T_6858;
  wire  _T_6859;
  wire [23:0] _T_6860;
  wire [24:0] _T_6861;
  wire [32:0] _T_6862;
  wire [33:0] _T_6863;
  wire [32:0] _T_6864;
  wire [31:0] _T_6866_number;
  wire [7:0] _T_6876;
  wire [7:0] _T_6878;
  wire [23:0] _T_6880;
  wire [7:0] _T_6881;
  wire [23:0] _T_6883;
  wire [31:0] _T_6884;
  wire [31:0] _T_6885;
  wire [31:0] _T_6894_number;
  wire [31:0] _T_6896_number;
  wire [31:0] _T_6904;
  wire [31:0] _T_6909_number;
  wire [31:0] _T_6919;
  wire  _T_6934;
  wire [32:0] _T_6936_number;
  wire [32:0] _T_6938_number;
  wire [7:0] _T_6944;
  wire [7:0] _T_6946;
  wire [24:0] _T_6948;
  wire [7:0] _T_6949;
  wire  _T_6950;
  wire [23:0] _T_6951;
  wire [24:0] _T_6952;
  wire [32:0] _T_6953;
  wire [33:0] _T_6967;
  wire [32:0] _T_6968;
  wire [31:0] _T_6970_number;
  wire [7:0] _T_6980;
  wire [7:0] _T_6982;
  wire [23:0] _T_6984;
  wire [7:0] _T_6985;
  wire [23:0] _T_6987;
  wire [31:0] _T_6988;
  wire [31:0] _T_6989;
  wire  RetimeWrapper_137_clock;
  wire  RetimeWrapper_137_reset;
  wire  RetimeWrapper_137_io_flow;
  wire  RetimeWrapper_137_io_in;
  wire  RetimeWrapper_137_io_out;
  wire  _T_6995;
  wire  _T_6997;
  wire  RetimeWrapper_138_clock;
  wire  RetimeWrapper_138_reset;
  wire  RetimeWrapper_138_io_flow;
  wire  RetimeWrapper_138_io_in;
  wire  RetimeWrapper_138_io_out;
  wire  _T_7002;
  wire  _T_7005;
  wire  _T_7008;
  wire  _T_7009;
  wire  _T_7010;
  wire [31:0] _T_7014;
  wire [63:0] _T_7015;
  wire [31:0] _T_7020_number;
  wire [31:0] _T_7022_number;
  wire [31:0] _T_7030;
  wire [31:0] _T_7035_number;
  wire [33:0] _GEN_2;
  wire [33:0] _T_7036;
  wire [5:0] x3244;
  wire [31:0] _T_7038_number;
  wire [33:0] _GEN_3;
  wire [33:0] _T_7039;
  wire [32:0] _T_7041_number;
  wire [32:0] _T_7043_number;
  wire [32:0] _T_7045_number;
  wire [32:0] _T_7053;
  wire  _T_7056;
  wire [32:0] _T_7058;
  wire [32:0] _T_7066;
  wire  _T_7069;
  wire [32:0] _T_7071;
  wire [33:0] _T_7072;
  wire [33:0] _T_7073;
  wire [32:0] _T_7074;
  wire [31:0] _T_7076_number;
  wire [31:0] _T_7090;
  wire [31:0] _T_7094;
  wire [32:0] _T_7096_number;
  wire [32:0] _T_7098_number;
  wire [32:0] _T_7100_number;
  wire [32:0] _T_7108;
  wire [32:0] _T_7121;
  wire  _T_7124;
  wire [32:0] _T_7126;
  wire [33:0] _T_7127;
  wire [32:0] _T_7128;
  wire [31:0] _T_7130_number;
  wire [31:0] _T_7144;
  wire [31:0] _T_7148;
  wire [5:0] x3251;
  wire [31:0] _T_7154_number;
  wire [31:0] _T_7164;
  wire  _T_7179;
  wire [32:0] _T_7185_number;
  wire [32:0] _T_7189_number;
  wire [32:0] _T_7210;
  wire  _T_7213;
  wire [32:0] _T_7215;
  wire [33:0] _T_7216;
  wire [33:0] _T_7217;
  wire [32:0] _T_7218;
  wire [31:0] _T_7220_number;
  wire [31:0] _T_7234;
  wire [31:0] _T_7238;
  wire [31:0] _T_7243;
  wire [31:0] _T_7245_number;
  wire [1:0] _T_7250;
  wire [29:0] _T_7251;
  wire [31:0] _T_7252;
  wire [31:0] _T_7254_number;
  wire  _T_7255;
  wire [1:0] _T_7259;
  wire [29:0] _T_7260;
  wire [31:0] _T_7261;
  wire [32:0] _T_7263_number;
  wire [32:0] _T_7265_number;
  wire [32:0] _T_7267_number;
  wire [32:0] _T_7275;
  wire  _T_7278;
  wire [32:0] _T_7280;
  wire [32:0] _T_7288;
  wire  _T_7291;
  wire [32:0] _T_7293;
  wire [33:0] _T_7294;
  wire [32:0] _T_7295;
  wire [31:0] _T_7297_number;
  wire [31:0] _T_7311;
  wire [31:0] _T_7315;
  wire [32:0] _T_7317_number;
  wire [32:0] _T_7319_number;
  wire [32:0] _T_7321_number;
  wire [32:0] _T_7329;
  wire [32:0] _T_7342;
  wire [33:0] _T_7348;
  wire [32:0] _T_7349;
  wire [31:0] _T_7351_number;
  wire [31:0] _T_7365;
  wire [31:0] _T_7369;
  wire [32:0] _T_7371_number;
  wire [32:0] _T_7373_number;
  wire [32:0] _T_7375_number;
  wire [32:0] _T_7383;
  wire  _T_7386;
  wire [32:0] _T_7388;
  wire [32:0] _T_7396;
  wire  _T_7399;
  wire [32:0] _T_7401;
  wire [33:0] _T_7402;
  wire [32:0] _T_7403;
  wire [31:0] _T_7405_number;
  wire [31:0] _T_7419;
  wire [31:0] _T_7423;
  wire [32:0] _T_7425_number;
  wire [32:0] _T_7427_number;
  wire [32:0] _T_7429_number;
  wire [32:0] _T_7437;
  wire [32:0] _T_7450;
  wire [33:0] _T_7456;
  wire [32:0] _T_7457;
  wire [31:0] _T_7459_number;
  wire [31:0] _T_7473;
  wire [31:0] _T_7477;
  wire [32:0] _T_7479_number;
  wire [32:0] _T_7481_number;
  wire [32:0] _T_7483_number;
  wire [32:0] _T_7491;
  wire  _T_7494;
  wire [32:0] _T_7496;
  wire [32:0] _T_7504;
  wire [32:0] _T_7509;
  wire [33:0] _T_7510;
  wire [32:0] _T_7511;
  wire [31:0] _T_7513_number;
  wire [31:0] _T_7527;
  wire [31:0] _T_7531;
  wire [63:0] _T_7539;
  wire  _T_7542;
  wire [31:0] _T_7546;
  wire [63:0] _T_7548;
  wire [63:0] _T_7550_number;
  wire [63:0] _T_7552_number;
  wire [63:0] _T_7560;
  wire [64:0] _T_7565_number;
  wire [64:0] _T_7567_number;
  wire [64:0] _T_7569_number;
  wire [64:0] _T_7577;
  wire  _T_7580;
  wire [64:0] _T_7582;
  wire [64:0] _T_7590;
  wire  _T_7593;
  wire [64:0] _T_7595;
  wire [65:0] _T_7596;
  wire [64:0] _T_7597;
  wire [63:0] _T_7599_number;
  wire [63:0] _T_7613;
  wire [63:0] _T_7617;
  wire [63:0] _T_7625;
  wire [32:0] _T_7630;
  wire [96:0] _T_7631;
  wire  _T_7637;
  wire  _T_7638;
  wire  _T_7645;
  wire [63:0] _T_7646;
  wire [95:0] _T_7647;
  wire [95:0] _T_7650_0;
  wire  _T_7664_0;
  wire [31:0] _T_7669_number;
  wire [31:0] _T_7671_number;
  wire [31:0] _T_7679;
  wire [31:0] _T_7684_number;
  wire [33:0] _GEN_4;
  wire [33:0] _T_7685;
  wire [5:0] x3371;
  wire [31:0] _T_7687_number;
  wire [33:0] _GEN_5;
  wire [33:0] _T_7688;
  wire [32:0] _T_7690_number;
  wire [32:0] _T_7692_number;
  wire [32:0] _T_7694_number;
  wire [32:0] _T_7702;
  wire  _T_7705;
  wire [32:0] _T_7707;
  wire [32:0] _T_7715;
  wire  _T_7718;
  wire [32:0] _T_7720;
  wire [33:0] _T_7721;
  wire [33:0] _T_7722;
  wire [32:0] _T_7723;
  wire [31:0] _T_7725_number;
  wire [31:0] _T_7739;
  wire [31:0] _T_7743;
  wire [32:0] _T_7745_number;
  wire [32:0] _T_7747_number;
  wire [32:0] _T_7749_number;
  wire [32:0] _T_7757;
  wire [32:0] _T_7770;
  wire  _T_7773;
  wire [32:0] _T_7775;
  wire [33:0] _T_7776;
  wire [32:0] _T_7777;
  wire [31:0] _T_7779_number;
  wire [31:0] _T_7793;
  wire [31:0] _T_7797;
  wire [5:0] x3378;
  wire [31:0] _T_7803_number;
  wire [31:0] _T_7813;
  wire  _T_7828;
  wire [32:0] _T_7834_number;
  wire [32:0] _T_7838_number;
  wire [32:0] _T_7859;
  wire  _T_7862;
  wire [32:0] _T_7864;
  wire [33:0] _T_7865;
  wire [33:0] _T_7866;
  wire [32:0] _T_7867;
  wire [31:0] _T_7869_number;
  wire [31:0] _T_7883;
  wire [31:0] _T_7887;
  wire [31:0] _T_7892;
  wire [31:0] _T_7894_number;
  wire [1:0] _T_7899;
  wire [29:0] _T_7900;
  wire [31:0] _T_7901;
  wire [31:0] _T_7903_number;
  wire  _T_7904;
  wire [1:0] _T_7908;
  wire [29:0] _T_7909;
  wire [31:0] _T_7910;
  wire [32:0] _T_7912_number;
  wire [32:0] _T_7914_number;
  wire [32:0] _T_7916_number;
  wire [32:0] _T_7924;
  wire  _T_7927;
  wire [32:0] _T_7929;
  wire [32:0] _T_7937;
  wire  _T_7940;
  wire [32:0] _T_7942;
  wire [33:0] _T_7943;
  wire [32:0] _T_7944;
  wire [31:0] _T_7946_number;
  wire [31:0] _T_7960;
  wire [31:0] _T_7964;
  wire [32:0] _T_7966_number;
  wire [32:0] _T_7968_number;
  wire [32:0] _T_7970_number;
  wire [32:0] _T_7978;
  wire [32:0] _T_7991;
  wire [33:0] _T_7997;
  wire [32:0] _T_7998;
  wire [31:0] _T_8000_number;
  wire [31:0] _T_8014;
  wire [31:0] _T_8018;
  wire [32:0] _T_8020_number;
  wire [32:0] _T_8022_number;
  wire [32:0] _T_8024_number;
  wire [32:0] _T_8032;
  wire  _T_8035;
  wire [32:0] _T_8037;
  wire [32:0] _T_8045;
  wire  _T_8048;
  wire [32:0] _T_8050;
  wire [33:0] _T_8051;
  wire [32:0] _T_8052;
  wire [31:0] _T_8054_number;
  wire [31:0] _T_8068;
  wire [31:0] _T_8072;
  wire [32:0] _T_8074_number;
  wire [32:0] _T_8076_number;
  wire [32:0] _T_8078_number;
  wire [32:0] _T_8086;
  wire [32:0] _T_8099;
  wire [33:0] _T_8105;
  wire [32:0] _T_8106;
  wire [31:0] _T_8108_number;
  wire [31:0] _T_8122;
  wire [31:0] _T_8126;
  wire [32:0] _T_8128_number;
  wire [32:0] _T_8130_number;
  wire [32:0] _T_8132_number;
  wire [32:0] _T_8140;
  wire  _T_8143;
  wire [32:0] _T_8145;
  wire [32:0] _T_8153;
  wire [32:0] _T_8158;
  wire [33:0] _T_8159;
  wire [32:0] _T_8160;
  wire [31:0] _T_8162_number;
  wire [31:0] _T_8176;
  wire [31:0] _T_8180;
  wire [63:0] _T_8188;
  wire  _T_8191;
  wire [31:0] _T_8195;
  wire [63:0] _T_8197;
  wire [63:0] _T_8199_number;
  wire [63:0] _T_8201_number;
  wire [63:0] _T_8209;
  wire [64:0] _T_8214_number;
  wire [64:0] _T_8216_number;
  wire [64:0] _T_8218_number;
  wire [64:0] _T_8226;
  wire  _T_8229;
  wire [64:0] _T_8231;
  wire [64:0] _T_8239;
  wire  _T_8242;
  wire [64:0] _T_8244;
  wire [65:0] _T_8245;
  wire [64:0] _T_8246;
  wire [63:0] _T_8248_number;
  wire [63:0] _T_8262;
  wire [63:0] _T_8266;
  wire [63:0] _T_8274;
  wire [32:0] _T_8279;
  wire [96:0] _T_8280;
  wire  _T_8286;
  wire  _T_8287;
  wire  _T_8294;
  wire [63:0] _T_8295;
  wire [95:0] _T_8296;
  wire [95:0] _T_8299_0;
  wire  _T_8313_0;
  wire  _T_8317;
  wire  _T_8320;
  wire  _T_8321;
  reg  _T_8324;
  reg [31:0] _RAND_17;
  wire  _T_8330;
  wire  _T_8333;
  wire  _T_8334;
  wire  _T_8335;
  wire  _T_8336;
  reg  _T_8339;
  reg [31:0] _RAND_18;
  wire  _T_8345;
  wire  RetimeWrapper_139_clock;
  wire  RetimeWrapper_139_reset;
  wire  RetimeWrapper_139_io_flow;
  wire  RetimeWrapper_139_io_in;
  wire  RetimeWrapper_139_io_out;
  wire  _T_8349;
  wire  _T_8351;
  wire  RetimeWrapper_140_clock;
  wire  RetimeWrapper_140_reset;
  wire  RetimeWrapper_140_io_flow;
  wire  RetimeWrapper_140_io_in;
  wire  RetimeWrapper_140_io_out;
  wire  _T_8357;
  wire  _T_8359;
  wire  _T_8363;
  wire  _T_8366;
  wire  _T_8367;
  reg  _T_8370;
  reg [31:0] _RAND_19;
  wire  _T_8376;
  wire  _T_8379;
  wire  _T_8380;
  wire  _T_8381;
  wire  _T_8382;
  reg  _T_8385;
  reg [31:0] _RAND_20;
  wire  _T_8391;
  wire  RetimeWrapper_141_clock;
  wire  RetimeWrapper_141_reset;
  wire  RetimeWrapper_141_io_flow;
  wire  RetimeWrapper_141_io_in;
  wire  RetimeWrapper_141_io_out;
  wire  _T_8395;
  wire  _T_8397;
  wire  RetimeWrapper_142_clock;
  wire  RetimeWrapper_142_reset;
  wire  RetimeWrapper_142_io_flow;
  wire  RetimeWrapper_142_io_in;
  wire  RetimeWrapper_142_io_out;
  wire  _T_8403;
  wire  _T_8405;
  wire [32:0] _T_8410_number;
  wire [32:0] _T_8412_number;
  wire [32:0] _T_8414_number;
  wire [32:0] _T_8422;
  wire  _T_8425;
  wire [32:0] _T_8427;
  wire [32:0] _T_8435;
  wire  _T_8438;
  wire [32:0] _T_8440;
  wire [33:0] _T_8441;
  wire [33:0] _T_8442;
  wire [32:0] _T_8443;
  wire [31:0] _T_8445_number;
  wire [31:0] _T_8459;
  wire [31:0] _T_8463;
  wire [31:0] _T_8471_number;
  wire [31:0] _T_8490;
  wire [31:0] _T_8495;
  wire  _T_8496;
  wire [31:0] _T_8501_number;
  wire  _T_8559;
  wire  _T_8560;
  wire  RetimeWrapper_143_clock;
  wire  RetimeWrapper_143_reset;
  wire  RetimeWrapper_143_io_flow;
  wire  RetimeWrapper_143_io_in;
  wire  RetimeWrapper_143_io_out;
  wire  _T_8564;
  wire  _T_8565;
  wire  _T_8566;
  wire  RetimeWrapper_144_clock;
  wire  RetimeWrapper_144_reset;
  wire  RetimeWrapper_144_io_flow;
  wire  RetimeWrapper_144_io_in;
  wire  RetimeWrapper_144_io_out;
  wire  _T_8571;
  wire  _T_8573;
  wire  RetimeWrapper_145_clock;
  wire  RetimeWrapper_145_reset;
  wire  RetimeWrapper_145_io_flow;
  wire  RetimeWrapper_145_io_in;
  wire  RetimeWrapper_145_io_out;
  wire  _T_8577;
  wire  _T_8579;
  wire  RetimeWrapper_146_clock;
  wire  RetimeWrapper_146_reset;
  wire  RetimeWrapper_146_io_flow;
  wire  RetimeWrapper_146_io_in;
  wire  RetimeWrapper_146_io_out;
  wire  _T_8583;
  wire  _T_8585;
  wire  RetimeWrapper_147_clock;
  wire  RetimeWrapper_147_reset;
  wire  RetimeWrapper_147_io_flow;
  wire  RetimeWrapper_147_io_in;
  wire  RetimeWrapper_147_io_out;
  wire  _T_8589;
  wire  _T_8591;
  wire  RetimeWrapper_148_clock;
  wire  RetimeWrapper_148_reset;
  wire  RetimeWrapper_148_io_flow;
  wire  RetimeWrapper_148_io_in;
  wire  RetimeWrapper_148_io_out;
  wire  _T_8595;
  wire  _T_8597;
  wire  RetimeWrapper_149_clock;
  wire  RetimeWrapper_149_reset;
  wire  RetimeWrapper_149_io_flow;
  wire  RetimeWrapper_149_io_in;
  wire  RetimeWrapper_149_io_out;
  wire  _T_8601;
  wire  _T_8603;
  wire  RetimeWrapper_150_clock;
  wire  RetimeWrapper_150_reset;
  wire  RetimeWrapper_150_io_flow;
  wire  RetimeWrapper_150_io_in;
  wire  RetimeWrapper_150_io_out;
  wire  _T_8607;
  wire  _T_8609;
  wire  RetimeWrapper_151_clock;
  wire  RetimeWrapper_151_reset;
  wire  RetimeWrapper_151_io_flow;
  wire  RetimeWrapper_151_io_in;
  wire  RetimeWrapper_151_io_out;
  wire  _T_8613;
  wire  _T_8615;
  wire  RetimeWrapper_152_clock;
  wire  RetimeWrapper_152_reset;
  wire  RetimeWrapper_152_io_flow;
  wire  RetimeWrapper_152_io_in;
  wire  RetimeWrapper_152_io_out;
  wire  _T_8619;
  wire  _T_8621;
  wire  RetimeWrapper_153_clock;
  wire  RetimeWrapper_153_reset;
  wire  RetimeWrapper_153_io_flow;
  wire  RetimeWrapper_153_io_in;
  wire  RetimeWrapper_153_io_out;
  wire  _T_8625;
  wire  _T_8627;
  wire  _T_8630;
  wire  _T_8633;
  wire  _T_8636;
  wire  _T_8639;
  wire  _T_8642;
  wire  RetimeWrapper_154_clock;
  wire  RetimeWrapper_154_reset;
  wire  RetimeWrapper_154_io_flow;
  wire  RetimeWrapper_154_io_in;
  wire  RetimeWrapper_154_io_out;
  wire  _T_8661;
  wire  _T_8663;
  wire  RetimeWrapper_155_clock;
  wire  RetimeWrapper_155_reset;
  wire  RetimeWrapper_155_io_flow;
  wire  RetimeWrapper_155_io_in;
  wire  RetimeWrapper_155_io_out;
  wire  _T_8667;
  wire  _T_8669;
  wire  RetimeWrapper_156_clock;
  wire  RetimeWrapper_156_reset;
  wire  RetimeWrapper_156_io_flow;
  wire  RetimeWrapper_156_io_in;
  wire  RetimeWrapper_156_io_out;
  wire  _T_8673;
  wire  _T_8675;
  wire  RetimeWrapper_157_clock;
  wire  RetimeWrapper_157_reset;
  wire  RetimeWrapper_157_io_flow;
  wire  RetimeWrapper_157_io_in;
  wire  RetimeWrapper_157_io_out;
  wire  _T_8679;
  wire  _T_8681;
  wire  RetimeWrapper_158_clock;
  wire  RetimeWrapper_158_reset;
  wire  RetimeWrapper_158_io_flow;
  wire  RetimeWrapper_158_io_in;
  wire  RetimeWrapper_158_io_out;
  wire  _T_8685;
  wire  _T_8687;
  wire  RetimeWrapper_159_clock;
  wire  RetimeWrapper_159_reset;
  wire  RetimeWrapper_159_io_flow;
  wire  RetimeWrapper_159_io_in;
  wire  RetimeWrapper_159_io_out;
  wire  _T_8691;
  wire  _T_8693;
  wire  RetimeWrapper_160_clock;
  wire  RetimeWrapper_160_reset;
  wire  RetimeWrapper_160_io_flow;
  wire  RetimeWrapper_160_io_in;
  wire  RetimeWrapper_160_io_out;
  wire  _T_8697;
  wire  _T_8699;
  wire  RetimeWrapper_161_clock;
  wire  RetimeWrapper_161_reset;
  wire  RetimeWrapper_161_io_flow;
  wire  RetimeWrapper_161_io_in;
  wire  RetimeWrapper_161_io_out;
  wire  _T_8703;
  wire  _T_8705;
  wire  RetimeWrapper_162_clock;
  wire  RetimeWrapper_162_reset;
  wire  RetimeWrapper_162_io_flow;
  wire  RetimeWrapper_162_io_in;
  wire  RetimeWrapper_162_io_out;
  wire  _T_8709;
  wire  _T_8711;
  wire  RetimeWrapper_163_clock;
  wire  RetimeWrapper_163_reset;
  wire  RetimeWrapper_163_io_flow;
  wire  RetimeWrapper_163_io_in;
  wire  RetimeWrapper_163_io_out;
  wire  _T_8715;
  wire  _T_8717;
  wire  RetimeWrapper_164_clock;
  wire  RetimeWrapper_164_reset;
  wire  RetimeWrapper_164_io_flow;
  wire  RetimeWrapper_164_io_in;
  wire  RetimeWrapper_164_io_out;
  wire  _T_8721;
  wire  _T_8723;
  wire  RetimeWrapper_165_clock;
  wire  RetimeWrapper_165_reset;
  wire  RetimeWrapper_165_io_flow;
  wire  RetimeWrapper_165_io_in;
  wire  RetimeWrapper_165_io_out;
  wire  _T_8727;
  wire  _T_8729;
  wire  RetimeWrapper_166_clock;
  wire  RetimeWrapper_166_reset;
  wire  RetimeWrapper_166_io_flow;
  wire  RetimeWrapper_166_io_in;
  wire  RetimeWrapper_166_io_out;
  wire  _T_8733;
  wire  _T_8735;
  wire  RetimeWrapper_167_clock;
  wire  RetimeWrapper_167_reset;
  wire  RetimeWrapper_167_io_flow;
  wire  RetimeWrapper_167_io_in;
  wire  RetimeWrapper_167_io_out;
  wire  _T_8739;
  wire  _T_8741;
  wire  RetimeWrapper_168_clock;
  wire  RetimeWrapper_168_reset;
  wire  RetimeWrapper_168_io_flow;
  wire  RetimeWrapper_168_io_in;
  wire  RetimeWrapper_168_io_out;
  wire  _T_8745;
  wire  _T_8747;
  wire  RetimeWrapper_169_clock;
  wire  RetimeWrapper_169_reset;
  wire  RetimeWrapper_169_io_flow;
  wire  RetimeWrapper_169_io_in;
  wire  RetimeWrapper_169_io_out;
  wire  _T_8751;
  wire  _T_8753;
  wire  RetimeWrapper_170_clock;
  wire  RetimeWrapper_170_reset;
  wire  RetimeWrapper_170_io_flow;
  wire  RetimeWrapper_170_io_in;
  wire  RetimeWrapper_170_io_out;
  wire  _T_8757;
  wire  _T_8759;
  wire  RetimeWrapper_171_clock;
  wire  RetimeWrapper_171_reset;
  wire  RetimeWrapper_171_io_flow;
  wire  RetimeWrapper_171_io_in;
  wire  RetimeWrapper_171_io_out;
  wire  _T_8763;
  wire  _T_8765;
  wire  RetimeWrapper_172_clock;
  wire  RetimeWrapper_172_reset;
  wire  RetimeWrapper_172_io_flow;
  wire  RetimeWrapper_172_io_in;
  wire  RetimeWrapper_172_io_out;
  wire  _T_8769;
  wire  _T_8771;
  wire  RetimeWrapper_173_clock;
  wire  RetimeWrapper_173_reset;
  wire  RetimeWrapper_173_io_flow;
  wire  RetimeWrapper_173_io_in;
  wire  RetimeWrapper_173_io_out;
  wire  _T_8775;
  wire  _T_8777;
  wire  RetimeWrapper_174_clock;
  wire  RetimeWrapper_174_reset;
  wire  RetimeWrapper_174_io_flow;
  wire  RetimeWrapper_174_io_in;
  wire  RetimeWrapper_174_io_out;
  wire  _T_8781;
  wire  _T_8783;
  wire  RetimeWrapper_175_clock;
  wire  RetimeWrapper_175_reset;
  wire  RetimeWrapper_175_io_flow;
  wire  RetimeWrapper_175_io_in;
  wire  RetimeWrapper_175_io_out;
  wire  _T_8787;
  wire  _T_8789;
  wire [31:0] _T_8790;
  wire [31:0] _T_8791;
  wire [31:0] _T_8792;
  wire [31:0] _T_8793;
  wire  _T_8794;
  wire  _T_8795;
  wire  _T_8796;
  wire  _T_8797;
  wire  _T_8800;
  wire  _T_8801;
  wire  _T_8805;
  wire  _T_8809;
  wire  _T_8813;
  wire [5:0] _T_8821_0_addr_0;
  wire  _T_8821_0_en;
  wire [5:0] _T_8821_1_addr_0;
  wire  _T_8821_1_en;
  wire [5:0] _T_8821_2_addr_0;
  wire  _T_8821_2_en;
  wire [5:0] _T_8821_3_addr_0;
  wire  _T_8821_3_en;
  wire [31:0] x3474_0_number;
  wire [31:0] x3474_1_number;
  wire [31:0] x3474_2_number;
  wire [31:0] x3474_3_number;
  wire [5:0] _T_8871_0_addr_0;
  wire  _T_8871_0_en;
  wire [5:0] _T_8871_1_addr_0;
  wire  _T_8871_1_en;
  wire [5:0] _T_8871_2_addr_0;
  wire  _T_8871_2_en;
  wire [5:0] _T_8871_3_addr_0;
  wire  _T_8871_3_en;
  wire [31:0] x3479_0_number;
  wire [31:0] x3479_1_number;
  wire [31:0] x3479_2_number;
  wire [31:0] x3479_3_number;
  wire [31:0] _T_8899_number;
  wire  _T_8900;
  wire [7:0] _T_8904;
  wire [39:0] _T_8905;
  wire  _T_8906;
  wire [7:0] _T_8910;
  wire [39:0] _T_8911;
  wire [79:0] _T_8912;
  wire [71:0] _T_8913;
  wire [31:0] _T_8915_number;
  wire [7:0] _T_8926;
  wire [7:0] _T_8928;
  wire [23:0] _T_8930;
  wire [7:0] _T_8931;
  wire [23:0] _T_8932;
  wire [31:0] _T_8933;
  wire [31:0] _T_8935_number;
  wire  _T_8936;
  wire [7:0] _T_8940;
  wire [39:0] _T_8941;
  wire  _T_8942;
  wire [7:0] _T_8946;
  wire [39:0] _T_8947;
  wire [79:0] _T_8948;
  wire [71:0] _T_8949;
  wire [31:0] _T_8951_number;
  wire [7:0] _T_8962;
  wire [7:0] _T_8964;
  wire [23:0] _T_8966;
  wire [7:0] _T_8967;
  wire [23:0] _T_8968;
  wire [31:0] _T_8969;
  wire [31:0] _T_8971_number;
  wire  _T_8972;
  wire [7:0] _T_8976;
  wire [39:0] _T_8977;
  wire  _T_8978;
  wire [7:0] _T_8982;
  wire [39:0] _T_8983;
  wire [79:0] _T_8984;
  wire [71:0] _T_8985;
  wire [31:0] _T_8987_number;
  wire [7:0] _T_8998;
  wire [7:0] _T_9000;
  wire [23:0] _T_9002;
  wire [7:0] _T_9003;
  wire [23:0] _T_9004;
  wire [31:0] _T_9005;
  wire [31:0] _T_9007_number;
  wire  _T_9008;
  wire [7:0] _T_9012;
  wire [39:0] _T_9013;
  wire  _T_9014;
  wire [7:0] _T_9018;
  wire [39:0] _T_9019;
  wire [79:0] _T_9020;
  wire [71:0] _T_9021;
  wire [31:0] _T_9023_number;
  wire [7:0] _T_9034;
  wire [7:0] _T_9036;
  wire [23:0] _T_9038;
  wire [7:0] _T_9039;
  wire [23:0] _T_9040;
  wire [31:0] _T_9041;
  wire [32:0] _T_9043_number;
  wire [32:0] _T_9045_number;
  wire [32:0] _T_9047_number;
  wire [7:0] _T_9051;
  wire [7:0] _T_9053;
  wire [24:0] _T_9055;
  wire [7:0] _T_9056;
  wire  _T_9057;
  wire [23:0] _T_9058;
  wire [24:0] _T_9059;
  wire [32:0] _T_9060;
  wire [7:0] _T_9064;
  wire [7:0] _T_9066;
  wire [24:0] _T_9068;
  wire [7:0] _T_9069;
  wire  _T_9070;
  wire [23:0] _T_9071;
  wire [24:0] _T_9072;
  wire [32:0] _T_9073;
  wire [33:0] _T_9074;
  wire [32:0] _T_9075;
  wire [31:0] _T_9077_number;
  wire [7:0] _T_9087;
  wire [7:0] _T_9089;
  wire [23:0] _T_9091;
  wire [7:0] _T_9092;
  wire [23:0] _T_9094;
  wire [31:0] _T_9095;
  wire [31:0] _T_9096;
  wire [32:0] _T_9099_number;
  wire [32:0] _T_9101_number;
  wire [32:0] _T_9103_number;
  wire [7:0] _T_9107;
  wire [7:0] _T_9109;
  wire [24:0] _T_9111;
  wire [7:0] _T_9112;
  wire  _T_9113;
  wire [23:0] _T_9114;
  wire [24:0] _T_9115;
  wire [32:0] _T_9116;
  wire [7:0] _T_9120;
  wire [7:0] _T_9122;
  wire [24:0] _T_9124;
  wire [7:0] _T_9125;
  wire  _T_9126;
  wire [23:0] _T_9127;
  wire [24:0] _T_9128;
  wire [32:0] _T_9129;
  wire [33:0] _T_9130;
  wire [32:0] _T_9131;
  wire [31:0] _T_9133_number;
  wire [7:0] _T_9143;
  wire [7:0] _T_9145;
  wire [23:0] _T_9147;
  wire [7:0] _T_9148;
  wire [23:0] _T_9150;
  wire [31:0] _T_9151;
  wire [31:0] _T_9152;
  wire  _T_9153;
  wire [32:0] _T_9155_number;
  wire [32:0] _T_9157_number;
  wire [32:0] _T_9159_number;
  wire [7:0] _T_9163;
  wire [7:0] _T_9165;
  wire [24:0] _T_9167;
  wire [7:0] _T_9168;
  wire  _T_9169;
  wire [23:0] _T_9170;
  wire [24:0] _T_9171;
  wire [32:0] _T_9172;
  wire [7:0] _T_9176;
  wire [7:0] _T_9178;
  wire [24:0] _T_9180;
  wire [7:0] _T_9181;
  wire  _T_9182;
  wire [23:0] _T_9183;
  wire [24:0] _T_9184;
  wire [32:0] _T_9185;
  wire [33:0] _T_9186;
  wire [32:0] _T_9187;
  wire [31:0] _T_9189_number;
  wire [7:0] _T_9199;
  wire [7:0] _T_9201;
  wire [23:0] _T_9203;
  wire [7:0] _T_9204;
  wire [23:0] _T_9206;
  wire [31:0] _T_9207;
  wire [31:0] _T_9208;
  wire [31:0] _T_9217_number;
  wire [31:0] _T_9227;
  wire  _T_9242;
  wire [32:0] _T_9244_number;
  wire [32:0] _T_9246_number;
  wire [7:0] _T_9252;
  wire [7:0] _T_9254;
  wire [24:0] _T_9256;
  wire [7:0] _T_9257;
  wire  _T_9258;
  wire [23:0] _T_9259;
  wire [24:0] _T_9260;
  wire [32:0] _T_9261;
  wire [33:0] _T_9275;
  wire [32:0] _T_9276;
  wire [31:0] _T_9278_number;
  wire [7:0] _T_9288;
  wire [7:0] _T_9290;
  wire [23:0] _T_9292;
  wire [7:0] _T_9293;
  wire [23:0] _T_9295;
  wire [31:0] _T_9296;
  wire [31:0] _T_9297;
  wire  _T_9300;
  wire  _T_9303;
  wire  _T_9304;
  wire  RetimeWrapper_176_clock;
  wire  RetimeWrapper_176_reset;
  wire  RetimeWrapper_176_io_flow;
  wire  RetimeWrapper_176_io_in;
  wire  RetimeWrapper_176_io_out;
  wire  _T_9309;
  wire  _T_9311;
  wire  _T_9312;
  wire  RetimeWrapper_177_clock;
  wire  RetimeWrapper_177_reset;
  wire  RetimeWrapper_177_io_flow;
  wire  RetimeWrapper_177_io_in;
  wire  RetimeWrapper_177_io_out;
  wire  _T_9316;
  wire  _T_9318;
  wire  _T_9320;
  wire  _T_9321;
  wire  _T_9324;
  wire  _T_9325;
  wire  _T_9326;
  wire  _T_9327;
  reg  _T_9330;
  reg [31:0] _RAND_21;
  wire  _T_9336;
  wire  RetimeWrapper_178_clock;
  wire  RetimeWrapper_178_reset;
  wire  RetimeWrapper_178_io_flow;
  wire  RetimeWrapper_178_io_in;
  wire  RetimeWrapper_178_io_out;
  wire  _T_9341;
  wire  _T_9343;
  wire  RetimeWrapper_179_clock;
  wire  RetimeWrapper_179_reset;
  wire  RetimeWrapper_179_io_flow;
  wire  RetimeWrapper_179_io_in;
  wire  RetimeWrapper_179_io_out;
  wire  _T_9350;
  wire  _T_9352;
  wire  _T_9359;
  wire [63:0] _T_9360;
  wire [31:0] _T_9361;
  wire  _T_9362;
  wire  _T_9363;
  wire  _T_9368;
  wire  _T_9369;
  wire  _T_9371;
  wire  RetimeWrapper_180_clock;
  wire  RetimeWrapper_180_reset;
  wire  RetimeWrapper_180_io_flow;
  wire  RetimeWrapper_180_io_in;
  wire  RetimeWrapper_180_io_out;
  wire  _T_9382;
  wire  _T_9384;
  wire  RetimeWrapper_181_clock;
  wire  RetimeWrapper_181_reset;
  wire  RetimeWrapper_181_io_flow;
  wire  RetimeWrapper_181_io_in;
  wire  RetimeWrapper_181_io_out;
  wire  _T_9390;
  wire  _T_9392;
  wire  _T_9393;
  wire  RetimeWrapper_182_clock;
  wire  RetimeWrapper_182_reset;
  wire  RetimeWrapper_182_io_flow;
  wire  RetimeWrapper_182_io_in;
  wire  RetimeWrapper_182_io_out;
  wire  _T_9397;
  wire  _T_9399;
  wire  _T_9400;
  wire  _T_9401;
  wire  RetimeWrapper_183_clock;
  wire  RetimeWrapper_183_reset;
  wire  RetimeWrapper_183_io_flow;
  wire  RetimeWrapper_183_io_in;
  wire  RetimeWrapper_183_io_out;
  wire  _T_9405;
  wire  _T_9407;
  wire  _T_9409;
  wire  _T_9410;
  wire  RetimeWrapper_184_clock;
  wire  RetimeWrapper_184_reset;
  wire  RetimeWrapper_184_io_flow;
  wire  RetimeWrapper_184_io_in;
  wire  RetimeWrapper_184_io_out;
  wire  _T_9414;
  wire  _T_9416;
  wire  RetimeWrapper_185_clock;
  wire  RetimeWrapper_185_reset;
  wire  RetimeWrapper_185_io_flow;
  wire  RetimeWrapper_185_io_in;
  wire  RetimeWrapper_185_io_out;
  wire  _T_9420;
  wire  _T_9422;
  wire  _T_9423;
  wire  RetimeWrapper_186_clock;
  wire  RetimeWrapper_186_reset;
  wire  RetimeWrapper_186_io_flow;
  wire  RetimeWrapper_186_io_in;
  wire  RetimeWrapper_186_io_out;
  wire  _T_9427;
  wire  _T_9429;
  wire  _T_9430;
  wire  _T_9431;
  wire  RetimeWrapper_187_clock;
  wire  RetimeWrapper_187_reset;
  wire  RetimeWrapper_187_io_flow;
  wire  RetimeWrapper_187_io_in;
  wire  RetimeWrapper_187_io_out;
  wire  _T_9438;
  wire  _T_9440;
  wire  _T_9443;
  wire  _T_9444;
  wire  _T_9445;
  wire  _T_9446;
  reg  _T_9449;
  reg [31:0] _RAND_22;
  wire  _T_9455;
  wire  RetimeWrapper_188_clock;
  wire  RetimeWrapper_188_reset;
  wire  RetimeWrapper_188_io_flow;
  wire  RetimeWrapper_188_io_in;
  wire  RetimeWrapper_188_io_out;
  wire  _T_9459;
  wire  _T_9461;
  wire  RetimeWrapper_189_clock;
  wire  RetimeWrapper_189_reset;
  wire  RetimeWrapper_189_io_flow;
  wire  RetimeWrapper_189_io_in;
  wire  RetimeWrapper_189_io_out;
  wire  _T_9467;
  wire  _T_9469;
  wire [31:0] _T_9473;
  wire  _T_9742;
  wire  _T_9744;
  wire  _T_9745;
  wire  _T_9746;
  wire  RetimeWrapper_190_clock;
  wire  RetimeWrapper_190_reset;
  wire  RetimeWrapper_190_io_flow;
  wire  RetimeWrapper_190_io_in;
  wire  RetimeWrapper_190_io_out;
  wire  _T_9753;
  wire  _T_9755;
  wire  RetimeWrapper_191_clock;
  wire  RetimeWrapper_191_reset;
  wire  RetimeWrapper_191_io_flow;
  wire  RetimeWrapper_191_io_in;
  wire  RetimeWrapper_191_io_out;
  wire  _T_9759;
  wire  _T_9761;
  wire [31:0] _T_9838_number;
  wire [31:0] _T_9840_number;
  wire [31:0] _T_9848;
  wire [31:0] _T_9859;
  wire [31:0] _T_9863;
  wire [31:0] _T_9864;
  wire  _T_9865;
  wire  RetimeWrapper_192_clock;
  wire  RetimeWrapper_192_reset;
  wire  RetimeWrapper_192_io_flow;
  wire  RetimeWrapper_192_io_in;
  wire  RetimeWrapper_192_io_out;
  wire  _T_9899;
  wire  _T_9901;
  wire [31:0] _T_9903_number;
  wire [31:0] _T_9913;
  wire  _T_9928;
  wire  _T_9929;
  wire [31:0] _T_9930;
  wire [31:0] _T_9932_number;
  wire [31:0] _T_9934_number;
  wire [31:0] _T_9942;
  wire [31:0] _T_9953;
  wire [31:0] _T_9957;
  wire [31:0] _T_9958;
  wire  _T_9959;
  wire [31:0] _T_9961_number;
  wire [31:0] _T_9963_number;
  wire [31:0] _T_9971;
  wire [31:0] _T_9982;
  wire [31:0] _T_9986;
  wire [31:0] _T_9987;
  wire  _T_9988;
  wire  _T_9989;
  wire [32:0] _T_9991_number;
  wire [32:0] _T_9993_number;
  wire [32:0] _T_9995_number;
  wire [32:0] _T_10003;
  wire  _T_10006;
  wire [32:0] _T_10008;
  wire [32:0] _T_10016;
  wire  _T_10019;
  wire [32:0] _T_10021;
  wire [33:0] _T_10022;
  wire [33:0] _T_10023;
  wire [32:0] _T_10024;
  wire [31:0] _T_10026_number;
  wire [31:0] _T_10040;
  wire [31:0] _T_10044;
  wire  _T_10045;
  wire  _T_10048;
  wire  _T_10049;
  wire  _T_10054;
  wire [31:0] _T_10055;
  wire [31:0] _T_10056;
  wire [31:0] _T_10057;
  wire [31:0] _T_10058;
  wire  _T_10059;
  wire  _T_10060;
  wire  _T_10061;
  wire  _T_10062;
  wire  _T_10065;
  wire  _T_10066;
  wire  _T_10070;
  wire  _T_10074;
  wire  _T_10078;
  wire [5:0] _T_10086_0_addr_0;
  wire  _T_10086_0_en;
  wire [5:0] _T_10086_1_addr_0;
  wire  _T_10086_1_en;
  wire [5:0] _T_10086_2_addr_0;
  wire  _T_10086_2_en;
  wire [5:0] _T_10086_3_addr_0;
  wire  _T_10086_3_en;
  wire [31:0] x3438_0_number;
  wire [31:0] x3438_1_number;
  wire [31:0] x3438_2_number;
  wire [31:0] x3438_3_number;
  wire [5:0] _T_10136_0_addr_0;
  wire  _T_10136_0_en;
  wire [5:0] _T_10136_1_addr_0;
  wire  _T_10136_1_en;
  wire [5:0] _T_10136_2_addr_0;
  wire  _T_10136_2_en;
  wire [5:0] _T_10136_3_addr_0;
  wire  _T_10136_3_en;
  wire [31:0] x3443_0_number;
  wire [31:0] x3443_1_number;
  wire [31:0] x3443_2_number;
  wire [31:0] x3443_3_number;
  wire [31:0] _T_10164_number;
  wire  _T_10165;
  wire [7:0] _T_10169;
  wire [39:0] _T_10170;
  wire  _T_10171;
  wire [7:0] _T_10175;
  wire [39:0] _T_10176;
  wire [79:0] _T_10177;
  wire [71:0] _T_10178;
  wire [31:0] _T_10180_number;
  wire [7:0] _T_10191;
  wire [7:0] _T_10193;
  wire [23:0] _T_10195;
  wire [7:0] _T_10196;
  wire [23:0] _T_10197;
  wire [31:0] _T_10198;
  wire [31:0] _T_10200_number;
  wire  _T_10201;
  wire [7:0] _T_10205;
  wire [39:0] _T_10206;
  wire  _T_10207;
  wire [7:0] _T_10211;
  wire [39:0] _T_10212;
  wire [79:0] _T_10213;
  wire [71:0] _T_10214;
  wire [31:0] _T_10216_number;
  wire [7:0] _T_10227;
  wire [7:0] _T_10229;
  wire [23:0] _T_10231;
  wire [7:0] _T_10232;
  wire [23:0] _T_10233;
  wire [31:0] _T_10234;
  wire [31:0] _T_10236_number;
  wire  _T_10237;
  wire [7:0] _T_10241;
  wire [39:0] _T_10242;
  wire  _T_10243;
  wire [7:0] _T_10247;
  wire [39:0] _T_10248;
  wire [79:0] _T_10249;
  wire [71:0] _T_10250;
  wire [31:0] _T_10252_number;
  wire [7:0] _T_10263;
  wire [7:0] _T_10265;
  wire [23:0] _T_10267;
  wire [7:0] _T_10268;
  wire [23:0] _T_10269;
  wire [31:0] _T_10270;
  wire [31:0] _T_10272_number;
  wire  _T_10273;
  wire [7:0] _T_10277;
  wire [39:0] _T_10278;
  wire  _T_10279;
  wire [7:0] _T_10283;
  wire [39:0] _T_10284;
  wire [79:0] _T_10285;
  wire [71:0] _T_10286;
  wire [31:0] _T_10288_number;
  wire [7:0] _T_10299;
  wire [7:0] _T_10301;
  wire [23:0] _T_10303;
  wire [7:0] _T_10304;
  wire [23:0] _T_10305;
  wire [31:0] _T_10306;
  wire [32:0] _T_10308_number;
  wire [32:0] _T_10310_number;
  wire [32:0] _T_10312_number;
  wire [7:0] _T_10316;
  wire [7:0] _T_10318;
  wire [24:0] _T_10320;
  wire [7:0] _T_10321;
  wire  _T_10322;
  wire [23:0] _T_10323;
  wire [24:0] _T_10324;
  wire [32:0] _T_10325;
  wire [7:0] _T_10329;
  wire [7:0] _T_10331;
  wire [24:0] _T_10333;
  wire [7:0] _T_10334;
  wire  _T_10335;
  wire [23:0] _T_10336;
  wire [24:0] _T_10337;
  wire [32:0] _T_10338;
  wire [33:0] _T_10339;
  wire [32:0] _T_10340;
  wire [31:0] _T_10342_number;
  wire [7:0] _T_10352;
  wire [7:0] _T_10354;
  wire [23:0] _T_10356;
  wire [7:0] _T_10357;
  wire [23:0] _T_10359;
  wire [31:0] _T_10360;
  wire [31:0] _T_10361;
  wire [32:0] _T_10364_number;
  wire [32:0] _T_10366_number;
  wire [32:0] _T_10368_number;
  wire [7:0] _T_10372;
  wire [7:0] _T_10374;
  wire [24:0] _T_10376;
  wire [7:0] _T_10377;
  wire  _T_10378;
  wire [23:0] _T_10379;
  wire [24:0] _T_10380;
  wire [32:0] _T_10381;
  wire [7:0] _T_10385;
  wire [7:0] _T_10387;
  wire [24:0] _T_10389;
  wire [7:0] _T_10390;
  wire  _T_10391;
  wire [23:0] _T_10392;
  wire [24:0] _T_10393;
  wire [32:0] _T_10394;
  wire [33:0] _T_10395;
  wire [32:0] _T_10396;
  wire [31:0] _T_10398_number;
  wire [7:0] _T_10408;
  wire [7:0] _T_10410;
  wire [23:0] _T_10412;
  wire [7:0] _T_10413;
  wire [23:0] _T_10415;
  wire [31:0] _T_10416;
  wire [31:0] _T_10417;
  wire  _T_10418;
  wire [32:0] _T_10420_number;
  wire [32:0] _T_10422_number;
  wire [32:0] _T_10424_number;
  wire [7:0] _T_10428;
  wire [7:0] _T_10430;
  wire [24:0] _T_10432;
  wire [7:0] _T_10433;
  wire  _T_10434;
  wire [23:0] _T_10435;
  wire [24:0] _T_10436;
  wire [32:0] _T_10437;
  wire [7:0] _T_10441;
  wire [7:0] _T_10443;
  wire [24:0] _T_10445;
  wire [7:0] _T_10446;
  wire  _T_10447;
  wire [23:0] _T_10448;
  wire [24:0] _T_10449;
  wire [32:0] _T_10450;
  wire [33:0] _T_10451;
  wire [32:0] _T_10452;
  wire [31:0] _T_10454_number;
  wire [7:0] _T_10464;
  wire [7:0] _T_10466;
  wire [23:0] _T_10468;
  wire [7:0] _T_10469;
  wire [23:0] _T_10471;
  wire [31:0] _T_10472;
  wire [31:0] _T_10473;
  wire [31:0] _T_10482_number;
  wire [31:0] _T_10492;
  wire  _T_10507;
  wire [32:0] _T_10509_number;
  wire [32:0] _T_10511_number;
  wire [7:0] _T_10517;
  wire [7:0] _T_10519;
  wire [24:0] _T_10521;
  wire [7:0] _T_10522;
  wire  _T_10523;
  wire [23:0] _T_10524;
  wire [24:0] _T_10525;
  wire [32:0] _T_10526;
  wire [33:0] _T_10540;
  wire [32:0] _T_10541;
  wire [31:0] _T_10543_number;
  wire [7:0] _T_10553;
  wire [7:0] _T_10555;
  wire [23:0] _T_10557;
  wire [7:0] _T_10558;
  wire [23:0] _T_10560;
  wire [31:0] _T_10561;
  wire [31:0] _T_10562;
  wire  _T_10565;
  wire  _T_10568;
  wire  _T_10569;
  wire  RetimeWrapper_193_clock;
  wire  RetimeWrapper_193_reset;
  wire  RetimeWrapper_193_io_flow;
  wire  RetimeWrapper_193_io_in;
  wire  RetimeWrapper_193_io_out;
  wire  _T_10574;
  wire  _T_10576;
  wire  _T_10577;
  wire  RetimeWrapper_194_clock;
  wire  RetimeWrapper_194_reset;
  wire  RetimeWrapper_194_io_flow;
  wire  RetimeWrapper_194_io_in;
  wire  RetimeWrapper_194_io_out;
  wire  _T_10581;
  wire [31:0] _T_10584_number;
  wire [31:0] _T_10586_number;
  wire [31:0] _T_10594;
  wire [31:0] _T_10599_number;
  wire [33:0] _GEN_6;
  wire [33:0] _T_10600;
  wire [5:0] x3308;
  wire [31:0] _T_10602_number;
  wire [33:0] _GEN_7;
  wire [33:0] _T_10603;
  wire [32:0] _T_10605_number;
  wire [32:0] _T_10607_number;
  wire [32:0] _T_10609_number;
  wire [32:0] _T_10617;
  wire  _T_10620;
  wire [32:0] _T_10622;
  wire [32:0] _T_10630;
  wire  _T_10633;
  wire [32:0] _T_10635;
  wire [33:0] _T_10636;
  wire [33:0] _T_10637;
  wire [32:0] _T_10638;
  wire [31:0] _T_10640_number;
  wire [31:0] _T_10654;
  wire [31:0] _T_10658;
  wire [32:0] _T_10660_number;
  wire [32:0] _T_10662_number;
  wire [32:0] _T_10664_number;
  wire [32:0] _T_10672;
  wire [32:0] _T_10685;
  wire  _T_10688;
  wire [32:0] _T_10690;
  wire [33:0] _T_10691;
  wire [32:0] _T_10692;
  wire [31:0] _T_10694_number;
  wire [31:0] _T_10708;
  wire [31:0] _T_10712;
  wire [5:0] x3315;
  wire [31:0] _T_10718_number;
  wire [31:0] _T_10728;
  wire  _T_10743;
  wire [32:0] _T_10749_number;
  wire [32:0] _T_10753_number;
  wire [32:0] _T_10774;
  wire  _T_10777;
  wire [32:0] _T_10779;
  wire [33:0] _T_10780;
  wire [33:0] _T_10781;
  wire [32:0] _T_10782;
  wire [31:0] _T_10784_number;
  wire [31:0] _T_10798;
  wire [31:0] _T_10802;
  wire [31:0] _T_10807;
  wire [31:0] _T_10809_number;
  wire [1:0] _T_10814;
  wire [29:0] _T_10815;
  wire [31:0] _T_10816;
  wire [31:0] _T_10818_number;
  wire  _T_10819;
  wire [1:0] _T_10823;
  wire [29:0] _T_10824;
  wire [31:0] _T_10825;
  wire [32:0] _T_10827_number;
  wire [32:0] _T_10829_number;
  wire [32:0] _T_10831_number;
  wire [32:0] _T_10839;
  wire  _T_10842;
  wire [32:0] _T_10844;
  wire [32:0] _T_10852;
  wire  _T_10855;
  wire [32:0] _T_10857;
  wire [33:0] _T_10858;
  wire [32:0] _T_10859;
  wire [31:0] _T_10861_number;
  wire [31:0] _T_10875;
  wire [31:0] _T_10879;
  wire [32:0] _T_10881_number;
  wire [32:0] _T_10883_number;
  wire [32:0] _T_10885_number;
  wire [32:0] _T_10893;
  wire [32:0] _T_10906;
  wire [33:0] _T_10912;
  wire [32:0] _T_10913;
  wire [31:0] _T_10915_number;
  wire [31:0] _T_10929;
  wire [31:0] _T_10933;
  wire [32:0] _T_10935_number;
  wire [32:0] _T_10937_number;
  wire [32:0] _T_10939_number;
  wire [32:0] _T_10947;
  wire  _T_10950;
  wire [32:0] _T_10952;
  wire [32:0] _T_10960;
  wire  _T_10963;
  wire [32:0] _T_10965;
  wire [33:0] _T_10966;
  wire [32:0] _T_10967;
  wire [31:0] _T_10969_number;
  wire [31:0] _T_10983;
  wire [31:0] _T_10987;
  wire [32:0] _T_10989_number;
  wire [32:0] _T_10991_number;
  wire [32:0] _T_10993_number;
  wire [32:0] _T_11001;
  wire [32:0] _T_11014;
  wire [33:0] _T_11020;
  wire [32:0] _T_11021;
  wire [31:0] _T_11023_number;
  wire [31:0] _T_11037;
  wire [31:0] _T_11041;
  wire [32:0] _T_11043_number;
  wire [32:0] _T_11045_number;
  wire [32:0] _T_11047_number;
  wire [32:0] _T_11055;
  wire  _T_11058;
  wire [32:0] _T_11060;
  wire [32:0] _T_11068;
  wire [32:0] _T_11073;
  wire [33:0] _T_11074;
  wire [32:0] _T_11075;
  wire [31:0] _T_11077_number;
  wire [31:0] _T_11091;
  wire [31:0] _T_11095;
  wire [63:0] _T_11103;
  wire  _T_11106;
  wire [31:0] _T_11110;
  wire [63:0] _T_11112;
  wire [63:0] _T_11114_number;
  wire [63:0] _T_11116_number;
  wire [63:0] _T_11124;
  wire [64:0] _T_11129_number;
  wire [64:0] _T_11131_number;
  wire [64:0] _T_11133_number;
  wire [64:0] _T_11141;
  wire  _T_11144;
  wire [64:0] _T_11146;
  wire [64:0] _T_11154;
  wire  _T_11157;
  wire [64:0] _T_11159;
  wire [65:0] _T_11160;
  wire [64:0] _T_11161;
  wire [63:0] _T_11163_number;
  wire [63:0] _T_11177;
  wire [63:0] _T_11181;
  wire [63:0] _T_11189;
  wire [32:0] _T_11194;
  wire [96:0] _T_11195;
  wire  _T_11201;
  wire  _T_11202;
  wire  _T_11209;
  wire [63:0] _T_11210;
  wire [95:0] _T_11211;
  wire [95:0] _T_11214_0;
  wire  _T_11228_0;
  wire [95:0] x3276;
  wire  _T_11238;
  wire  _T_11239;
  wire  _T_11240;
  wire  _T_11243_0;
  wire [95:0] _T_11250_0;
  wire [31:0] _T_11254;
  wire  _T_11259;
  wire  RetimeWrapper_195_clock;
  wire  RetimeWrapper_195_reset;
  wire  RetimeWrapper_195_io_flow;
  wire  RetimeWrapper_195_io_in;
  wire  RetimeWrapper_195_io_out;
  wire  _T_11263;
  wire  _T_11264;
  wire  _T_11265;
  wire [31:0] _T_11266;
  wire  RetimeWrapper_196_clock;
  wire  RetimeWrapper_196_reset;
  wire  RetimeWrapper_196_io_flow;
  wire  RetimeWrapper_196_io_in;
  wire  RetimeWrapper_196_io_out;
  wire  _T_11275;
  wire  _T_11277;
  wire [31:0] _T_11278;
  wire  RetimeWrapper_197_clock;
  wire  RetimeWrapper_197_reset;
  wire  RetimeWrapper_197_io_flow;
  wire  RetimeWrapper_197_io_in;
  wire  RetimeWrapper_197_io_out;
  wire  _T_11287;
  wire  _T_11289;
  wire [32:0] _T_11291_number;
  wire [32:0] _T_11293_number;
  wire [32:0] _T_11295_number;
  wire [32:0] _T_11303;
  wire  _T_11306;
  wire [32:0] _T_11308;
  wire [32:0] _T_11316;
  wire  _T_11319;
  wire [32:0] _T_11321;
  wire [33:0] _T_11322;
  wire [33:0] _T_11323;
  wire [32:0] _T_11324;
  wire [31:0] _T_11326_number;
  wire [31:0] _T_11340;
  wire [31:0] _T_11344;
  wire [31:0] _T_11352_number;
  wire [31:0] _T_11371;
  wire [31:0] _T_11376;
  wire  _T_11377;
  wire [31:0] _T_11382_number;
  wire  _T_11440;
  wire  _T_11441;
  wire  RetimeWrapper_198_clock;
  wire  RetimeWrapper_198_reset;
  wire  RetimeWrapper_198_io_flow;
  wire  RetimeWrapper_198_io_in;
  wire  RetimeWrapper_198_io_out;
  wire  _T_11445;
  wire  _T_11446;
  wire  _T_11447;
  wire  _T_11449;
  wire  _T_11451;
  wire  _T_11454;
  wire  _T_11455;
  wire  _T_11456;
  wire  _T_11457;
  reg  _T_11460;
  reg [31:0] _RAND_23;
  wire  _T_11466;
  wire  RetimeWrapper_199_clock;
  wire  RetimeWrapper_199_reset;
  wire  RetimeWrapper_199_io_flow;
  wire  RetimeWrapper_199_io_in;
  wire  RetimeWrapper_199_io_out;
  wire  _T_11470;
  wire  _T_11472;
  wire  RetimeWrapper_200_clock;
  wire  RetimeWrapper_200_reset;
  wire  RetimeWrapper_200_io_flow;
  wire  RetimeWrapper_200_io_in;
  wire  RetimeWrapper_200_io_out;
  wire  _T_11478;
  wire  _T_11480;
  wire [31:0] _T_11484;
  wire  _T_11753;
  wire  _T_11755;
  wire  _T_11756;
  wire  _T_11757;
  wire  RetimeWrapper_201_clock;
  wire  RetimeWrapper_201_reset;
  wire  RetimeWrapper_201_io_flow;
  wire  RetimeWrapper_201_io_in;
  wire  RetimeWrapper_201_io_out;
  wire  _T_11764;
  wire  _T_11766;
  wire  RetimeWrapper_202_clock;
  wire  RetimeWrapper_202_reset;
  wire  RetimeWrapper_202_io_flow;
  wire  RetimeWrapper_202_io_in;
  wire  RetimeWrapper_202_io_out;
  wire  _T_11770;
  wire  _T_11772;
  wire [31:0] _T_11849_number;
  wire [31:0] _T_11851_number;
  wire [31:0] _T_11859;
  wire [31:0] _T_11870;
  wire [31:0] _T_11874;
  wire [31:0] _T_11875;
  wire  _T_11876;
  wire  RetimeWrapper_203_clock;
  wire  RetimeWrapper_203_reset;
  wire  RetimeWrapper_203_io_flow;
  wire  RetimeWrapper_203_io_in;
  wire  RetimeWrapper_203_io_out;
  wire  _T_11910;
  wire  _T_11912;
  wire [31:0] _T_11914_number;
  wire [31:0] _T_11924;
  wire  _T_11939;
  wire  _T_11940;
  wire [31:0] _T_11941;
  wire [31:0] _T_11943_number;
  wire [31:0] _T_11945_number;
  wire [31:0] _T_11953;
  wire [31:0] _T_11964;
  wire [31:0] _T_11968;
  wire [31:0] _T_11969;
  wire  _T_11970;
  wire [31:0] _T_11972_number;
  wire [31:0] _T_11974_number;
  wire [31:0] _T_11982;
  wire [31:0] _T_11993;
  wire [31:0] _T_11997;
  wire [31:0] _T_11998;
  wire  _T_11999;
  wire  _T_12000;
  wire [32:0] _T_12002_number;
  wire [32:0] _T_12004_number;
  wire [32:0] _T_12006_number;
  wire [32:0] _T_12014;
  wire  _T_12017;
  wire [32:0] _T_12019;
  wire [32:0] _T_12027;
  wire  _T_12030;
  wire [32:0] _T_12032;
  wire [33:0] _T_12033;
  wire [33:0] _T_12034;
  wire [32:0] _T_12035;
  wire [31:0] _T_12037_number;
  wire [31:0] _T_12051;
  wire [31:0] _T_12055;
  wire  _T_12056;
  wire  _T_12059;
  wire  _T_12060;
  wire  _T_12065;
  wire [95:0] x3213;
  wire  _T_12072;
  wire  _T_12073;
  wire  _T_12074;
  wire  _T_12077_0;
  wire [95:0] _T_12084_0;
  wire [31:0] _T_12088;
  wire  _T_12093;
  wire  RetimeWrapper_204_clock;
  wire  RetimeWrapper_204_reset;
  wire  RetimeWrapper_204_io_flow;
  wire  RetimeWrapper_204_io_in;
  wire  RetimeWrapper_204_io_out;
  wire  _T_12097;
  wire  _T_12098;
  wire  _T_12099;
  wire [31:0] _T_12100;
  wire  RetimeWrapper_205_clock;
  wire  RetimeWrapper_205_reset;
  wire  RetimeWrapper_205_io_flow;
  wire  RetimeWrapper_205_io_in;
  wire  RetimeWrapper_205_io_out;
  wire  _T_12109;
  wire  _T_12111;
  wire [31:0] _T_12112;
  wire  RetimeWrapper_206_clock;
  wire  RetimeWrapper_206_reset;
  wire  RetimeWrapper_206_io_flow;
  wire  RetimeWrapper_206_io_in;
  wire  RetimeWrapper_206_io_out;
  wire  _T_12121;
  wire  _T_12123;
  wire [31:0] _T_12124;
  wire [31:0] _T_12126_number;
  wire [31:0] _T_12128_number;
  wire [31:0] _T_12136;
  wire [31:0] _T_12147;
  wire [31:0] _T_12151;
  wire [31:0] _T_12152;
  wire  _T_12153;
  wire [31:0] _T_12155_number;
  wire [31:0] _T_12157_number;
  wire [31:0] _T_12165;
  wire [31:0] _T_12176;
  wire [31:0] _T_12180;
  wire [31:0] _T_12181;
  wire  _T_12182;
  wire  _T_12183;
  wire [32:0] _T_12185_number;
  wire [32:0] _T_12187_number;
  wire [32:0] _T_12189_number;
  wire [32:0] _T_12197;
  wire  _T_12200;
  wire [32:0] _T_12202;
  wire [32:0] _T_12210;
  wire  _T_12213;
  wire [32:0] _T_12215;
  wire [33:0] _T_12216;
  wire [33:0] _T_12217;
  wire [32:0] _T_12218;
  wire [31:0] _T_12220_number;
  wire [31:0] _T_12234;
  wire [31:0] _T_12238;
  wire  _T_12239;
  wire  _T_12242;
  wire  _T_12243;
  wire  _T_12248;
  wire [31:0] _T_12249;
  wire [31:0] _T_12251_number;
  wire [31:0] _T_12253_number;
  wire [31:0] _T_12261;
  wire [31:0] _T_12272;
  wire [31:0] _T_12276;
  wire [31:0] _T_12277;
  wire  _T_12278;
  wire [31:0] _T_12280_number;
  wire [31:0] _T_12282_number;
  wire [31:0] _T_12290;
  wire [31:0] _T_12301;
  wire [31:0] _T_12305;
  wire [31:0] _T_12306;
  wire  _T_12307;
  wire  _T_12308;
  wire [32:0] _T_12310_number;
  wire [32:0] _T_12312_number;
  wire [32:0] _T_12314_number;
  wire [32:0] _T_12322;
  wire  _T_12325;
  wire [32:0] _T_12327;
  wire [32:0] _T_12335;
  wire  _T_12338;
  wire [32:0] _T_12340;
  wire [33:0] _T_12341;
  wire [33:0] _T_12342;
  wire [32:0] _T_12343;
  wire [31:0] _T_12345_number;
  wire [31:0] _T_12359;
  wire [31:0] _T_12363;
  wire  _T_12364;
  wire  _T_12367;
  wire  _T_12368;
  wire  _T_12373;
  wire [95:0] x3340;
  wire  _T_12380;
  wire  _T_12381;
  wire  _T_12382;
  wire  _T_12385_0;
  wire [95:0] _T_12392_0;
  wire [31:0] _T_12396;
  wire  _T_12401;
  wire  RetimeWrapper_207_clock;
  wire  RetimeWrapper_207_reset;
  wire  RetimeWrapper_207_io_flow;
  wire  RetimeWrapper_207_io_in;
  wire  RetimeWrapper_207_io_out;
  wire  _T_12405;
  wire  _T_12406;
  wire  _T_12407;
  wire [31:0] _T_12408;
  wire  RetimeWrapper_208_clock;
  wire  RetimeWrapper_208_reset;
  wire  RetimeWrapper_208_io_flow;
  wire  RetimeWrapper_208_io_in;
  wire  RetimeWrapper_208_io_out;
  wire  _T_12417;
  wire  _T_12419;
  wire [31:0] _T_12420;
  wire  RetimeWrapper_209_clock;
  wire  RetimeWrapper_209_reset;
  wire  RetimeWrapper_209_io_flow;
  wire  RetimeWrapper_209_io_in;
  wire  RetimeWrapper_209_io_out;
  wire  _T_12429;
  wire  _T_12431;
  wire [95:0] x3403;
  wire  _T_12438;
  wire  _T_12439;
  wire  _T_12440;
  wire  _T_12443_0;
  wire [95:0] _T_12450_0;
  wire [31:0] _T_12454;
  wire  _T_12459;
  wire  RetimeWrapper_210_clock;
  wire  RetimeWrapper_210_reset;
  wire  RetimeWrapper_210_io_flow;
  wire  RetimeWrapper_210_io_in;
  wire  RetimeWrapper_210_io_out;
  wire  _T_12463;
  wire  _T_12464;
  wire  _T_12465;
  wire [31:0] _T_12466;
  wire  RetimeWrapper_211_clock;
  wire  RetimeWrapper_211_reset;
  wire  RetimeWrapper_211_io_flow;
  wire  RetimeWrapper_211_io_in;
  wire  RetimeWrapper_211_io_out;
  wire  _T_12475;
  wire  _T_12477;
  wire [31:0] _T_12478;
  wire  RetimeWrapper_212_clock;
  wire  RetimeWrapper_212_reset;
  wire  RetimeWrapper_212_io_flow;
  wire  RetimeWrapper_212_io_in;
  wire  RetimeWrapper_212_io_out;
  wire  _T_12487;
  wire  _T_12489;
  RetimeWrapper RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  Seqpipe RootController_sm (
    .clock(RootController_sm_clock),
    .reset(RootController_sm_reset),
    .io_input_enable(RootController_sm_io_input_enable),
    .io_input_stageDone_0(RootController_sm_io_input_stageDone_0),
    .io_input_stageDone_1(RootController_sm_io_input_stageDone_1),
    .io_input_stageMask_0(RootController_sm_io_input_stageMask_0),
    .io_input_stageMask_1(RootController_sm_io_input_stageMask_1),
    .io_input_rst(RootController_sm_io_input_rst),
    .io_output_done(RootController_sm_io_output_done),
    .io_output_stageEnable_0(RootController_sm_io_output_stageEnable_0),
    .io_output_stageEnable_1(RootController_sm_io_output_stageEnable_1),
    .io_output_rst_en(RootController_sm_io_output_rst_en)
  );
  FF_1 x3152_0 (
    .clock(x3152_0_clock),
    .reset(x3152_0_reset),
    .io_input_0_data(x3152_0_io_input_0_data),
    .io_input_0_init(x3152_0_io_input_0_init),
    .io_input_0_enable(x3152_0_io_input_0_enable),
    .io_input_0_reset(x3152_0_io_input_0_reset),
    .io_output_data(x3152_0_io_output_data)
  );
  SpecialAccum x3152_1 (
    .clock(x3152_1_clock),
    .reset(x3152_1_reset),
    .io_input_next(x3152_1_io_input_next),
    .io_input_enable(x3152_1_io_input_enable),
    .io_input_reset(x3152_1_io_input_reset),
    .io_output(x3152_1_io_output)
  );
  Counter x3155 (
    .clock(x3155_clock),
    .reset(x3155_reset),
    .io_input_stops_0(x3155_io_input_stops_0),
    .io_input_reset(x3155_io_input_reset),
    .io_input_enable(x3155_io_input_enable),
    .io_output_counts_1(x3155_io_output_counts_1),
    .io_output_counts_0(x3155_io_output_counts_0)
  );
  Metapipe x3515_sm (
    .clock(x3515_sm_clock),
    .reset(x3515_sm_reset),
    .io_input_enable(x3515_sm_io_input_enable),
    .io_input_numIter(x3515_sm_io_input_numIter),
    .io_input_stageDone_0(x3515_sm_io_input_stageDone_0),
    .io_input_stageDone_1(x3515_sm_io_input_stageDone_1),
    .io_input_stageDone_2(x3515_sm_io_input_stageDone_2),
    .io_input_stageDone_3(x3515_sm_io_input_stageDone_3),
    .io_input_stageDone_4(x3515_sm_io_input_stageDone_4),
    .io_input_rst(x3515_sm_io_input_rst),
    .io_output_done(x3515_sm_io_output_done),
    .io_output_stageEnable_0(x3515_sm_io_output_stageEnable_0),
    .io_output_stageEnable_1(x3515_sm_io_output_stageEnable_1),
    .io_output_stageEnable_2(x3515_sm_io_output_stageEnable_2),
    .io_output_stageEnable_3(x3515_sm_io_output_stageEnable_3),
    .io_output_stageEnable_4(x3515_sm_io_output_stageEnable_4),
    .io_output_rst_en(x3515_sm_io_output_rst_en),
    .io_output_ctr_inc(x3515_sm_io_output_ctr_inc)
  );
  NBufFF b1202_chain (
    .clock(b1202_chain_clock),
    .reset(b1202_chain_reset),
    .io_sEn_0(b1202_chain_io_sEn_0),
    .io_sEn_1(b1202_chain_io_sEn_1),
    .io_sEn_2(b1202_chain_io_sEn_2),
    .io_sEn_3(b1202_chain_io_sEn_3),
    .io_sEn_4(b1202_chain_io_sEn_4),
    .io_sDone_0(b1202_chain_io_sDone_0),
    .io_sDone_1(b1202_chain_io_sDone_1),
    .io_sDone_2(b1202_chain_io_sDone_2),
    .io_sDone_3(b1202_chain_io_sDone_3),
    .io_sDone_4(b1202_chain_io_sDone_4),
    .io_input_0_data(b1202_chain_io_input_0_data),
    .io_input_0_enable(b1202_chain_io_input_0_enable),
    .io_input_0_reset(b1202_chain_io_input_0_reset),
    .io_output_1_data(b1202_chain_io_output_1_data),
    .io_output_2_data(b1202_chain_io_output_2_data),
    .io_output_4_data(b1202_chain_io_output_4_data)
  );
  NBufFF b1203_chain (
    .clock(b1203_chain_clock),
    .reset(b1203_chain_reset),
    .io_sEn_0(b1203_chain_io_sEn_0),
    .io_sEn_1(b1203_chain_io_sEn_1),
    .io_sEn_2(b1203_chain_io_sEn_2),
    .io_sEn_3(b1203_chain_io_sEn_3),
    .io_sEn_4(b1203_chain_io_sEn_4),
    .io_sDone_0(b1203_chain_io_sDone_0),
    .io_sDone_1(b1203_chain_io_sDone_1),
    .io_sDone_2(b1203_chain_io_sDone_2),
    .io_sDone_3(b1203_chain_io_sDone_3),
    .io_sDone_4(b1203_chain_io_sDone_4),
    .io_input_0_data(b1203_chain_io_input_0_data),
    .io_input_0_enable(b1203_chain_io_input_0_enable),
    .io_input_0_reset(b1203_chain_io_input_0_reset),
    .io_output_1_data(b1203_chain_io_output_1_data),
    .io_output_2_data(b1203_chain_io_output_2_data),
    .io_output_4_data(b1203_chain_io_output_4_data)
  );
  NBufFF_2 x3156_0 (
    .clock(x3156_0_clock),
    .reset(x3156_0_reset),
    .io_sEn_0(x3156_0_io_sEn_0),
    .io_sEn_1(x3156_0_io_sEn_1),
    .io_sEn_2(x3156_0_io_sEn_2),
    .io_sEn_3(x3156_0_io_sEn_3),
    .io_sDone_0(x3156_0_io_sDone_0),
    .io_sDone_1(x3156_0_io_sDone_1),
    .io_sDone_2(x3156_0_io_sDone_2),
    .io_sDone_3(x3156_0_io_sDone_3),
    .io_input_0_data(x3156_0_io_input_0_data),
    .io_input_0_enable(x3156_0_io_input_0_enable),
    .io_input_0_reset(x3156_0_io_input_0_reset),
    .io_output_1_data(x3156_0_io_output_1_data),
    .io_output_2_data(x3156_0_io_output_2_data),
    .io_output_3_data(x3156_0_io_output_3_data)
  );
  NBufFF_2 x3157_0 (
    .clock(x3157_0_clock),
    .reset(x3157_0_reset),
    .io_sEn_0(x3157_0_io_sEn_0),
    .io_sEn_1(x3157_0_io_sEn_1),
    .io_sEn_2(x3157_0_io_sEn_2),
    .io_sEn_3(x3157_0_io_sEn_3),
    .io_sDone_0(x3157_0_io_sDone_0),
    .io_sDone_1(x3157_0_io_sDone_1),
    .io_sDone_2(x3157_0_io_sDone_2),
    .io_sDone_3(x3157_0_io_sDone_3),
    .io_input_0_data(x3157_0_io_input_0_data),
    .io_input_0_enable(x3157_0_io_input_0_enable),
    .io_input_0_reset(x3157_0_io_input_0_reset),
    .io_output_1_data(x3157_0_io_output_1_data),
    .io_output_2_data(x3157_0_io_output_2_data),
    .io_output_3_data(x3157_0_io_output_3_data)
  );
  NBufSRAMnoBcast x3158_0 (
    .clock(x3158_0_clock),
    .reset(x3158_0_reset),
    .io_sEn_0(x3158_0_io_sEn_0),
    .io_sEn_1(x3158_0_io_sEn_1),
    .io_sEn_2(x3158_0_io_sEn_2),
    .io_sDone_0(x3158_0_io_sDone_0),
    .io_sDone_1(x3158_0_io_sDone_1),
    .io_sDone_2(x3158_0_io_sDone_2),
    .io_w_0_addr_0(x3158_0_io_w_0_addr_0),
    .io_w_0_data(x3158_0_io_w_0_data),
    .io_w_0_en(x3158_0_io_w_0_en),
    .io_r_0_addr_0(x3158_0_io_r_0_addr_0),
    .io_r_0_en(x3158_0_io_r_0_en),
    .io_r_1_addr_0(x3158_0_io_r_1_addr_0),
    .io_r_1_en(x3158_0_io_r_1_en),
    .io_r_2_addr_0(x3158_0_io_r_2_addr_0),
    .io_r_2_en(x3158_0_io_r_2_en),
    .io_r_3_addr_0(x3158_0_io_r_3_addr_0),
    .io_r_3_en(x3158_0_io_r_3_en),
    .io_output_data_8(x3158_0_io_output_data_8),
    .io_output_data_9(x3158_0_io_output_data_9),
    .io_output_data_10(x3158_0_io_output_data_10),
    .io_output_data_11(x3158_0_io_output_data_11)
  );
  NBufSRAMnoBcast x3159_0 (
    .clock(x3159_0_clock),
    .reset(x3159_0_reset),
    .io_sEn_0(x3159_0_io_sEn_0),
    .io_sEn_1(x3159_0_io_sEn_1),
    .io_sEn_2(x3159_0_io_sEn_2),
    .io_sDone_0(x3159_0_io_sDone_0),
    .io_sDone_1(x3159_0_io_sDone_1),
    .io_sDone_2(x3159_0_io_sDone_2),
    .io_w_0_addr_0(x3159_0_io_w_0_addr_0),
    .io_w_0_data(x3159_0_io_w_0_data),
    .io_w_0_en(x3159_0_io_w_0_en),
    .io_r_0_addr_0(x3159_0_io_r_0_addr_0),
    .io_r_0_en(x3159_0_io_r_0_en),
    .io_r_1_addr_0(x3159_0_io_r_1_addr_0),
    .io_r_1_en(x3159_0_io_r_1_en),
    .io_r_2_addr_0(x3159_0_io_r_2_addr_0),
    .io_r_2_en(x3159_0_io_r_2_en),
    .io_r_3_addr_0(x3159_0_io_r_3_addr_0),
    .io_r_3_en(x3159_0_io_r_3_en),
    .io_output_data_8(x3159_0_io_output_data_8),
    .io_output_data_9(x3159_0_io_output_data_9),
    .io_output_data_10(x3159_0_io_output_data_10),
    .io_output_data_11(x3159_0_io_output_data_11)
  );
  NBufSRAMnoBcast_2 x3160_0 (
    .clock(x3160_0_clock),
    .reset(x3160_0_reset),
    .io_sEn_0(x3160_0_io_sEn_0),
    .io_sEn_1(x3160_0_io_sEn_1),
    .io_sDone_0(x3160_0_io_sDone_0),
    .io_sDone_1(x3160_0_io_sDone_1),
    .io_w_0_addr_0(x3160_0_io_w_0_addr_0),
    .io_w_0_data(x3160_0_io_w_0_data),
    .io_w_0_en(x3160_0_io_w_0_en),
    .io_r_0_addr_0(x3160_0_io_r_0_addr_0),
    .io_r_0_en(x3160_0_io_r_0_en),
    .io_r_1_addr_0(x3160_0_io_r_1_addr_0),
    .io_r_1_en(x3160_0_io_r_1_en),
    .io_r_2_addr_0(x3160_0_io_r_2_addr_0),
    .io_r_2_en(x3160_0_io_r_2_en),
    .io_r_3_addr_0(x3160_0_io_r_3_addr_0),
    .io_r_3_en(x3160_0_io_r_3_en),
    .io_output_data_4(x3160_0_io_output_data_4),
    .io_output_data_5(x3160_0_io_output_data_5),
    .io_output_data_6(x3160_0_io_output_data_6),
    .io_output_data_7(x3160_0_io_output_data_7)
  );
  NBufSRAMnoBcast_2 x3161_0 (
    .clock(x3161_0_clock),
    .reset(x3161_0_reset),
    .io_sEn_0(x3161_0_io_sEn_0),
    .io_sEn_1(x3161_0_io_sEn_1),
    .io_sDone_0(x3161_0_io_sDone_0),
    .io_sDone_1(x3161_0_io_sDone_1),
    .io_w_0_addr_0(x3161_0_io_w_0_addr_0),
    .io_w_0_data(x3161_0_io_w_0_data),
    .io_w_0_en(x3161_0_io_w_0_en),
    .io_r_0_addr_0(x3161_0_io_r_0_addr_0),
    .io_r_0_en(x3161_0_io_r_0_en),
    .io_r_1_addr_0(x3161_0_io_r_1_addr_0),
    .io_r_1_en(x3161_0_io_r_1_en),
    .io_r_2_addr_0(x3161_0_io_r_2_addr_0),
    .io_r_2_en(x3161_0_io_r_2_en),
    .io_r_3_addr_0(x3161_0_io_r_3_addr_0),
    .io_r_3_en(x3161_0_io_r_3_en),
    .io_output_data_4(x3161_0_io_output_data_4),
    .io_output_data_5(x3161_0_io_output_data_5),
    .io_output_data_6(x3161_0_io_output_data_6),
    .io_output_data_7(x3161_0_io_output_data_7)
  );
  Parallel x3174_sm (
    .clock(x3174_sm_clock),
    .reset(x3174_sm_reset),
    .io_input_enable(x3174_sm_io_input_enable),
    .io_input_stageDone_0(x3174_sm_io_input_stageDone_0),
    .io_input_stageDone_1(x3174_sm_io_input_stageDone_1),
    .io_input_stageMask_0(x3174_sm_io_input_stageMask_0),
    .io_input_stageMask_1(x3174_sm_io_input_stageMask_1),
    .io_input_rst(x3174_sm_io_input_rst),
    .io_output_done(x3174_sm_io_output_done),
    .io_output_stageEnable_0(x3174_sm_io_output_stageEnable_0),
    .io_output_stageEnable_1(x3174_sm_io_output_stageEnable_1),
    .io_output_rst_en(x3174_sm_io_output_rst_en)
  );
  Innerpipe x3167_sm (
    .clock(x3167_sm_clock),
    .reset(x3167_sm_reset),
    .io_input_enable(x3167_sm_io_input_enable),
    .io_input_ctr_done(x3167_sm_io_input_ctr_done),
    .io_input_rst(x3167_sm_io_input_rst),
    .io_output_done(x3167_sm_io_output_done),
    .io_output_ctr_inc(x3167_sm_io_output_ctr_inc)
  );
  Innerpipe x3173_sm (
    .clock(x3173_sm_clock),
    .reset(x3173_sm_reset),
    .io_input_enable(x3173_sm_io_input_enable),
    .io_input_ctr_done(x3173_sm_io_input_ctr_done),
    .io_input_rst(x3173_sm_io_input_rst),
    .io_output_done(x3173_sm_io_output_done),
    .io_output_ctr_inc(x3173_sm_io_output_ctr_inc)
  );
  Parallel x3301_sm (
    .clock(x3301_sm_clock),
    .reset(x3301_sm_reset),
    .io_input_enable(x3301_sm_io_input_enable),
    .io_input_stageDone_0(x3301_sm_io_input_stageDone_0),
    .io_input_stageDone_1(x3301_sm_io_input_stageDone_1),
    .io_input_stageMask_0(x3301_sm_io_input_stageMask_0),
    .io_input_stageMask_1(x3301_sm_io_input_stageMask_1),
    .io_input_rst(x3301_sm_io_input_rst),
    .io_output_done(x3301_sm_io_output_done),
    .io_output_stageEnable_0(x3301_sm_io_output_stageEnable_0),
    .io_output_stageEnable_1(x3301_sm_io_output_stageEnable_1),
    .io_output_rst_en(x3301_sm_io_output_rst_en)
  );
  Parallel x3237_sm (
    .clock(x3237_sm_clock),
    .reset(x3237_sm_reset),
    .io_input_enable(x3237_sm_io_input_enable),
    .io_input_stageDone_0(x3237_sm_io_input_stageDone_0),
    .io_input_stageDone_1(x3237_sm_io_input_stageDone_1),
    .io_input_stageMask_0(x3237_sm_io_input_stageMask_0),
    .io_input_stageMask_1(x3237_sm_io_input_stageMask_1),
    .io_input_rst(x3237_sm_io_input_rst),
    .io_output_done(x3237_sm_io_output_done),
    .io_output_stageEnable_0(x3237_sm_io_output_stageEnable_0),
    .io_output_stageEnable_1(x3237_sm_io_output_stageEnable_1),
    .io_output_rst_en(x3237_sm_io_output_rst_en)
  );
  SRFF x3175_valid_srff (
    .clock(x3175_valid_srff_clock),
    .reset(x3175_valid_srff_reset),
    .io_input_set(x3175_valid_srff_io_input_set),
    .io_input_reset(x3175_valid_srff_io_input_reset),
    .io_input_asyn_reset(x3175_valid_srff_io_input_asyn_reset),
    .io_output_data(x3175_valid_srff_io_output_data)
  );
  GeneralFIFO x3176 (
    .clock(x3176_clock),
    .reset(x3176_reset),
    .io_in_0_data(x3176_io_in_0_data),
    .io_in_0_en(x3176_io_in_0_en),
    .io_out_0(x3176_io_out_0),
    .io_deq_0(x3176_io_deq_0),
    .io_empty(x3176_io_empty),
    .io_full(x3176_io_full)
  );
  Innerpipe x3208_sm (
    .clock(x3208_sm_clock),
    .reset(x3208_sm_reset),
    .io_input_enable(x3208_sm_io_input_enable),
    .io_input_ctr_done(x3208_sm_io_input_ctr_done),
    .io_input_rst(x3208_sm_io_input_rst),
    .io_output_done(x3208_sm_io_output_done),
    .io_output_ctr_inc(x3208_sm_io_output_ctr_inc)
  );
  Seqpipe x3236_sm (
    .clock(x3236_sm_clock),
    .reset(x3236_sm_reset),
    .io_input_enable(x3236_sm_io_input_enable),
    .io_input_stageDone_0(x3236_sm_io_input_stageDone_0),
    .io_input_stageDone_1(x3236_sm_io_input_stageDone_1),
    .io_input_stageMask_0(x3236_sm_io_input_stageMask_0),
    .io_input_stageMask_1(x3236_sm_io_input_stageMask_1),
    .io_input_rst(x3236_sm_io_input_rst),
    .io_output_done(x3236_sm_io_output_done),
    .io_output_stageEnable_0(x3236_sm_io_output_stageEnable_0),
    .io_output_stageEnable_1(x3236_sm_io_output_stageEnable_1),
    .io_output_rst_en(x3236_sm_io_output_rst_en)
  );
  FF_1 x3210_0 (
    .clock(x3210_0_clock),
    .reset(x3210_0_reset),
    .io_input_0_data(x3210_0_io_input_0_data),
    .io_input_0_init(x3210_0_io_input_0_init),
    .io_input_0_enable(x3210_0_io_input_0_enable),
    .io_input_0_reset(x3210_0_io_input_0_reset),
    .io_output_data(x3210_0_io_output_data)
  );
  FF_1 x3211_0 (
    .clock(x3211_0_clock),
    .reset(x3211_0_reset),
    .io_input_0_data(x3211_0_io_input_0_data),
    .io_input_0_init(x3211_0_io_input_0_init),
    .io_input_0_enable(x3211_0_io_input_0_enable),
    .io_input_0_reset(x3211_0_io_input_0_reset),
    .io_output_data(x3211_0_io_output_data)
  );
  FF_1 x3212_0 (
    .clock(x3212_0_clock),
    .reset(x3212_0_reset),
    .io_input_0_data(x3212_0_io_input_0_data),
    .io_input_0_init(x3212_0_io_input_0_init),
    .io_input_0_enable(x3212_0_io_input_0_enable),
    .io_input_0_reset(x3212_0_io_input_0_reset),
    .io_output_data(x3212_0_io_output_data)
  );
  Innerpipe x3220_sm (
    .clock(x3220_sm_clock),
    .reset(x3220_sm_reset),
    .io_input_enable(x3220_sm_io_input_enable),
    .io_input_ctr_done(x3220_sm_io_input_ctr_done),
    .io_input_rst(x3220_sm_io_input_rst),
    .io_output_done(x3220_sm_io_output_done),
    .io_output_ctr_inc(x3220_sm_io_output_ctr_inc)
  );
  Counter_1 x3223 (
    .clock(x3223_clock),
    .reset(x3223_reset),
    .io_input_stops_0(x3223_io_input_stops_0),
    .io_input_reset(x3223_io_input_reset),
    .io_input_enable(x3223_io_input_enable),
    .io_output_counts_0(x3223_io_output_counts_0),
    .io_output_done(x3223_io_output_done)
  );
  Streaminner x3235_sm (
    .io_input_ctr_done(x3235_sm_io_input_ctr_done),
    .io_output_done(x3235_sm_io_output_done)
  );
  Parallel x3300_sm (
    .clock(x3300_sm_clock),
    .reset(x3300_sm_reset),
    .io_input_enable(x3300_sm_io_input_enable),
    .io_input_stageDone_0(x3300_sm_io_input_stageDone_0),
    .io_input_stageDone_1(x3300_sm_io_input_stageDone_1),
    .io_input_stageMask_0(x3300_sm_io_input_stageMask_0),
    .io_input_stageMask_1(x3300_sm_io_input_stageMask_1),
    .io_input_rst(x3300_sm_io_input_rst),
    .io_output_done(x3300_sm_io_output_done),
    .io_output_stageEnable_0(x3300_sm_io_output_stageEnable_0),
    .io_output_stageEnable_1(x3300_sm_io_output_stageEnable_1),
    .io_output_rst_en(x3300_sm_io_output_rst_en)
  );
  SRFF x3238_valid_srff (
    .clock(x3238_valid_srff_clock),
    .reset(x3238_valid_srff_reset),
    .io_input_set(x3238_valid_srff_io_input_set),
    .io_input_reset(x3238_valid_srff_io_input_reset),
    .io_input_asyn_reset(x3238_valid_srff_io_input_asyn_reset),
    .io_output_data(x3238_valid_srff_io_output_data)
  );
  GeneralFIFO x3239 (
    .clock(x3239_clock),
    .reset(x3239_reset),
    .io_in_0_data(x3239_io_in_0_data),
    .io_in_0_en(x3239_io_in_0_en),
    .io_out_0(x3239_io_out_0),
    .io_deq_0(x3239_io_deq_0),
    .io_empty(x3239_io_empty),
    .io_full(x3239_io_full)
  );
  Innerpipe x3271_sm (
    .clock(x3271_sm_clock),
    .reset(x3271_sm_reset),
    .io_input_enable(x3271_sm_io_input_enable),
    .io_input_ctr_done(x3271_sm_io_input_ctr_done),
    .io_input_rst(x3271_sm_io_input_rst),
    .io_output_done(x3271_sm_io_output_done),
    .io_output_ctr_inc(x3271_sm_io_output_ctr_inc)
  );
  Seqpipe x3299_sm (
    .clock(x3299_sm_clock),
    .reset(x3299_sm_reset),
    .io_input_enable(x3299_sm_io_input_enable),
    .io_input_stageDone_0(x3299_sm_io_input_stageDone_0),
    .io_input_stageDone_1(x3299_sm_io_input_stageDone_1),
    .io_input_stageMask_0(x3299_sm_io_input_stageMask_0),
    .io_input_stageMask_1(x3299_sm_io_input_stageMask_1),
    .io_input_rst(x3299_sm_io_input_rst),
    .io_output_done(x3299_sm_io_output_done),
    .io_output_stageEnable_0(x3299_sm_io_output_stageEnable_0),
    .io_output_stageEnable_1(x3299_sm_io_output_stageEnable_1),
    .io_output_rst_en(x3299_sm_io_output_rst_en)
  );
  FF_1 x3273_0 (
    .clock(x3273_0_clock),
    .reset(x3273_0_reset),
    .io_input_0_data(x3273_0_io_input_0_data),
    .io_input_0_init(x3273_0_io_input_0_init),
    .io_input_0_enable(x3273_0_io_input_0_enable),
    .io_input_0_reset(x3273_0_io_input_0_reset),
    .io_output_data(x3273_0_io_output_data)
  );
  FF_1 x3274_0 (
    .clock(x3274_0_clock),
    .reset(x3274_0_reset),
    .io_input_0_data(x3274_0_io_input_0_data),
    .io_input_0_init(x3274_0_io_input_0_init),
    .io_input_0_enable(x3274_0_io_input_0_enable),
    .io_input_0_reset(x3274_0_io_input_0_reset),
    .io_output_data(x3274_0_io_output_data)
  );
  FF_1 x3275_0 (
    .clock(x3275_0_clock),
    .reset(x3275_0_reset),
    .io_input_0_data(x3275_0_io_input_0_data),
    .io_input_0_init(x3275_0_io_input_0_init),
    .io_input_0_enable(x3275_0_io_input_0_enable),
    .io_input_0_reset(x3275_0_io_input_0_reset),
    .io_output_data(x3275_0_io_output_data)
  );
  Innerpipe x3283_sm (
    .clock(x3283_sm_clock),
    .reset(x3283_sm_reset),
    .io_input_enable(x3283_sm_io_input_enable),
    .io_input_ctr_done(x3283_sm_io_input_ctr_done),
    .io_input_rst(x3283_sm_io_input_rst),
    .io_output_done(x3283_sm_io_output_done),
    .io_output_ctr_inc(x3283_sm_io_output_ctr_inc)
  );
  Counter_1 x3286 (
    .clock(x3286_clock),
    .reset(x3286_reset),
    .io_input_stops_0(x3286_io_input_stops_0),
    .io_input_reset(x3286_io_input_reset),
    .io_input_enable(x3286_io_input_enable),
    .io_output_counts_0(x3286_io_output_counts_0),
    .io_output_done(x3286_io_output_done)
  );
  Streaminner x3298_sm (
    .io_input_ctr_done(x3298_sm_io_input_ctr_done),
    .io_output_done(x3298_sm_io_output_done)
  );
  Parallel x3428_sm (
    .clock(x3428_sm_clock),
    .reset(x3428_sm_reset),
    .io_input_enable(x3428_sm_io_input_enable),
    .io_input_stageDone_0(x3428_sm_io_input_stageDone_0),
    .io_input_stageDone_1(x3428_sm_io_input_stageDone_1),
    .io_input_stageMask_0(x3428_sm_io_input_stageMask_0),
    .io_input_stageMask_1(x3428_sm_io_input_stageMask_1),
    .io_input_rst(x3428_sm_io_input_rst),
    .io_output_done(x3428_sm_io_output_done),
    .io_output_stageEnable_0(x3428_sm_io_output_stageEnable_0),
    .io_output_stageEnable_1(x3428_sm_io_output_stageEnable_1),
    .io_output_rst_en(x3428_sm_io_output_rst_en)
  );
  Parallel x3364_sm (
    .clock(x3364_sm_clock),
    .reset(x3364_sm_reset),
    .io_input_enable(x3364_sm_io_input_enable),
    .io_input_stageDone_0(x3364_sm_io_input_stageDone_0),
    .io_input_stageDone_1(x3364_sm_io_input_stageDone_1),
    .io_input_stageMask_0(x3364_sm_io_input_stageMask_0),
    .io_input_stageMask_1(x3364_sm_io_input_stageMask_1),
    .io_input_rst(x3364_sm_io_input_rst),
    .io_output_done(x3364_sm_io_output_done),
    .io_output_stageEnable_0(x3364_sm_io_output_stageEnable_0),
    .io_output_stageEnable_1(x3364_sm_io_output_stageEnable_1),
    .io_output_rst_en(x3364_sm_io_output_rst_en)
  );
  SRFF x3302_valid_srff (
    .clock(x3302_valid_srff_clock),
    .reset(x3302_valid_srff_reset),
    .io_input_set(x3302_valid_srff_io_input_set),
    .io_input_reset(x3302_valid_srff_io_input_reset),
    .io_input_asyn_reset(x3302_valid_srff_io_input_asyn_reset),
    .io_output_data(x3302_valid_srff_io_output_data)
  );
  GeneralFIFO x3303 (
    .clock(x3303_clock),
    .reset(x3303_reset),
    .io_in_0_data(x3303_io_in_0_data),
    .io_in_0_en(x3303_io_in_0_en),
    .io_out_0(x3303_io_out_0),
    .io_deq_0(x3303_io_deq_0),
    .io_empty(x3303_io_empty),
    .io_full(x3303_io_full)
  );
  Innerpipe x3335_sm (
    .clock(x3335_sm_clock),
    .reset(x3335_sm_reset),
    .io_input_enable(x3335_sm_io_input_enable),
    .io_input_ctr_done(x3335_sm_io_input_ctr_done),
    .io_input_rst(x3335_sm_io_input_rst),
    .io_output_done(x3335_sm_io_output_done),
    .io_output_ctr_inc(x3335_sm_io_output_ctr_inc)
  );
  Seqpipe x3363_sm (
    .clock(x3363_sm_clock),
    .reset(x3363_sm_reset),
    .io_input_enable(x3363_sm_io_input_enable),
    .io_input_stageDone_0(x3363_sm_io_input_stageDone_0),
    .io_input_stageDone_1(x3363_sm_io_input_stageDone_1),
    .io_input_stageMask_0(x3363_sm_io_input_stageMask_0),
    .io_input_stageMask_1(x3363_sm_io_input_stageMask_1),
    .io_input_rst(x3363_sm_io_input_rst),
    .io_output_done(x3363_sm_io_output_done),
    .io_output_stageEnable_0(x3363_sm_io_output_stageEnable_0),
    .io_output_stageEnable_1(x3363_sm_io_output_stageEnable_1),
    .io_output_rst_en(x3363_sm_io_output_rst_en)
  );
  FF_1 x3337_0 (
    .clock(x3337_0_clock),
    .reset(x3337_0_reset),
    .io_input_0_data(x3337_0_io_input_0_data),
    .io_input_0_init(x3337_0_io_input_0_init),
    .io_input_0_enable(x3337_0_io_input_0_enable),
    .io_input_0_reset(x3337_0_io_input_0_reset),
    .io_output_data(x3337_0_io_output_data)
  );
  FF_1 x3338_0 (
    .clock(x3338_0_clock),
    .reset(x3338_0_reset),
    .io_input_0_data(x3338_0_io_input_0_data),
    .io_input_0_init(x3338_0_io_input_0_init),
    .io_input_0_enable(x3338_0_io_input_0_enable),
    .io_input_0_reset(x3338_0_io_input_0_reset),
    .io_output_data(x3338_0_io_output_data)
  );
  FF_1 x3339_0 (
    .clock(x3339_0_clock),
    .reset(x3339_0_reset),
    .io_input_0_data(x3339_0_io_input_0_data),
    .io_input_0_init(x3339_0_io_input_0_init),
    .io_input_0_enable(x3339_0_io_input_0_enable),
    .io_input_0_reset(x3339_0_io_input_0_reset),
    .io_output_data(x3339_0_io_output_data)
  );
  Innerpipe x3347_sm (
    .clock(x3347_sm_clock),
    .reset(x3347_sm_reset),
    .io_input_enable(x3347_sm_io_input_enable),
    .io_input_ctr_done(x3347_sm_io_input_ctr_done),
    .io_input_rst(x3347_sm_io_input_rst),
    .io_output_done(x3347_sm_io_output_done),
    .io_output_ctr_inc(x3347_sm_io_output_ctr_inc)
  );
  Counter_1 x3350 (
    .clock(x3350_clock),
    .reset(x3350_reset),
    .io_input_stops_0(x3350_io_input_stops_0),
    .io_input_reset(x3350_io_input_reset),
    .io_input_enable(x3350_io_input_enable),
    .io_output_counts_0(x3350_io_output_counts_0),
    .io_output_done(x3350_io_output_done)
  );
  Streaminner x3362_sm (
    .io_input_ctr_done(x3362_sm_io_input_ctr_done),
    .io_output_done(x3362_sm_io_output_done)
  );
  Parallel x3427_sm (
    .clock(x3427_sm_clock),
    .reset(x3427_sm_reset),
    .io_input_enable(x3427_sm_io_input_enable),
    .io_input_stageDone_0(x3427_sm_io_input_stageDone_0),
    .io_input_stageDone_1(x3427_sm_io_input_stageDone_1),
    .io_input_stageMask_0(x3427_sm_io_input_stageMask_0),
    .io_input_stageMask_1(x3427_sm_io_input_stageMask_1),
    .io_input_rst(x3427_sm_io_input_rst),
    .io_output_done(x3427_sm_io_output_done),
    .io_output_stageEnable_0(x3427_sm_io_output_stageEnable_0),
    .io_output_stageEnable_1(x3427_sm_io_output_stageEnable_1),
    .io_output_rst_en(x3427_sm_io_output_rst_en)
  );
  SRFF x3365_valid_srff (
    .clock(x3365_valid_srff_clock),
    .reset(x3365_valid_srff_reset),
    .io_input_set(x3365_valid_srff_io_input_set),
    .io_input_reset(x3365_valid_srff_io_input_reset),
    .io_input_asyn_reset(x3365_valid_srff_io_input_asyn_reset),
    .io_output_data(x3365_valid_srff_io_output_data)
  );
  GeneralFIFO x3366 (
    .clock(x3366_clock),
    .reset(x3366_reset),
    .io_in_0_data(x3366_io_in_0_data),
    .io_in_0_en(x3366_io_in_0_en),
    .io_out_0(x3366_io_out_0),
    .io_deq_0(x3366_io_deq_0),
    .io_empty(x3366_io_empty),
    .io_full(x3366_io_full)
  );
  Innerpipe x3398_sm (
    .clock(x3398_sm_clock),
    .reset(x3398_sm_reset),
    .io_input_enable(x3398_sm_io_input_enable),
    .io_input_ctr_done(x3398_sm_io_input_ctr_done),
    .io_input_rst(x3398_sm_io_input_rst),
    .io_output_done(x3398_sm_io_output_done),
    .io_output_ctr_inc(x3398_sm_io_output_ctr_inc)
  );
  Seqpipe x3426_sm (
    .clock(x3426_sm_clock),
    .reset(x3426_sm_reset),
    .io_input_enable(x3426_sm_io_input_enable),
    .io_input_stageDone_0(x3426_sm_io_input_stageDone_0),
    .io_input_stageDone_1(x3426_sm_io_input_stageDone_1),
    .io_input_stageMask_0(x3426_sm_io_input_stageMask_0),
    .io_input_stageMask_1(x3426_sm_io_input_stageMask_1),
    .io_input_rst(x3426_sm_io_input_rst),
    .io_output_done(x3426_sm_io_output_done),
    .io_output_stageEnable_0(x3426_sm_io_output_stageEnable_0),
    .io_output_stageEnable_1(x3426_sm_io_output_stageEnable_1),
    .io_output_rst_en(x3426_sm_io_output_rst_en)
  );
  FF_1 x3400_0 (
    .clock(x3400_0_clock),
    .reset(x3400_0_reset),
    .io_input_0_data(x3400_0_io_input_0_data),
    .io_input_0_init(x3400_0_io_input_0_init),
    .io_input_0_enable(x3400_0_io_input_0_enable),
    .io_input_0_reset(x3400_0_io_input_0_reset),
    .io_output_data(x3400_0_io_output_data)
  );
  FF_1 x3401_0 (
    .clock(x3401_0_clock),
    .reset(x3401_0_reset),
    .io_input_0_data(x3401_0_io_input_0_data),
    .io_input_0_init(x3401_0_io_input_0_init),
    .io_input_0_enable(x3401_0_io_input_0_enable),
    .io_input_0_reset(x3401_0_io_input_0_reset),
    .io_output_data(x3401_0_io_output_data)
  );
  FF_1 x3402_0 (
    .clock(x3402_0_clock),
    .reset(x3402_0_reset),
    .io_input_0_data(x3402_0_io_input_0_data),
    .io_input_0_init(x3402_0_io_input_0_init),
    .io_input_0_enable(x3402_0_io_input_0_enable),
    .io_input_0_reset(x3402_0_io_input_0_reset),
    .io_output_data(x3402_0_io_output_data)
  );
  Innerpipe x3410_sm (
    .clock(x3410_sm_clock),
    .reset(x3410_sm_reset),
    .io_input_enable(x3410_sm_io_input_enable),
    .io_input_ctr_done(x3410_sm_io_input_ctr_done),
    .io_input_rst(x3410_sm_io_input_rst),
    .io_output_done(x3410_sm_io_output_done),
    .io_output_ctr_inc(x3410_sm_io_output_ctr_inc)
  );
  Counter_1 x3413 (
    .clock(x3413_clock),
    .reset(x3413_reset),
    .io_input_stops_0(x3413_io_input_stops_0),
    .io_input_reset(x3413_io_input_reset),
    .io_input_enable(x3413_io_input_enable),
    .io_output_counts_0(x3413_io_output_counts_0),
    .io_output_done(x3413_io_output_done)
  );
  Streaminner x3425_sm (
    .io_input_ctr_done(x3425_sm_io_input_ctr_done),
    .io_output_done(x3425_sm_io_output_done)
  );
  SpecialAccum x3429_0 (
    .clock(x3429_0_clock),
    .reset(x3429_0_reset),
    .io_input_next(x3429_0_io_input_next),
    .io_input_enable(x3429_0_io_input_enable),
    .io_input_reset(x3429_0_io_input_reset),
    .io_output(x3429_0_io_output)
  );
  NBufFF_4 x3429_1 (
    .clock(x3429_1_clock),
    .reset(x3429_1_reset),
    .io_sEn_0(x3429_1_io_sEn_0),
    .io_sEn_1(x3429_1_io_sEn_1),
    .io_sDone_0(x3429_1_io_sDone_0),
    .io_sDone_1(x3429_1_io_sDone_1),
    .io_input_0_data(x3429_1_io_input_0_data),
    .io_input_0_enable(x3429_1_io_input_0_enable),
    .io_input_0_reset(x3429_1_io_input_0_reset),
    .io_output_1_data(x3429_1_io_output_1_data)
  );
  SpecialAccum x3430_0 (
    .clock(x3430_0_clock),
    .reset(x3430_0_reset),
    .io_input_next(x3430_0_io_input_next),
    .io_input_enable(x3430_0_io_input_enable),
    .io_input_reset(x3430_0_io_input_reset),
    .io_output(x3430_0_io_output)
  );
  NBufFF_4 x3430_1 (
    .clock(x3430_1_clock),
    .reset(x3430_1_reset),
    .io_sEn_0(x3430_1_io_sEn_0),
    .io_sEn_1(x3430_1_io_sEn_1),
    .io_sDone_0(x3430_1_io_sDone_0),
    .io_sDone_1(x3430_1_io_sDone_1),
    .io_input_0_data(x3430_1_io_input_0_data),
    .io_input_0_enable(x3430_1_io_input_0_enable),
    .io_input_0_reset(x3430_1_io_input_0_reset),
    .io_output_1_data(x3430_1_io_output_1_data)
  );
  Parallel x3503_sm (
    .clock(x3503_sm_clock),
    .reset(x3503_sm_reset),
    .io_input_enable(x3503_sm_io_input_enable),
    .io_input_stageDone_0(x3503_sm_io_input_stageDone_0),
    .io_input_stageDone_1(x3503_sm_io_input_stageDone_1),
    .io_input_stageMask_0(x3503_sm_io_input_stageMask_0),
    .io_input_stageMask_1(x3503_sm_io_input_stageMask_1),
    .io_input_rst(x3503_sm_io_input_rst),
    .io_output_done(x3503_sm_io_output_done),
    .io_output_stageEnable_0(x3503_sm_io_output_stageEnable_0),
    .io_output_stageEnable_1(x3503_sm_io_output_stageEnable_1),
    .io_output_rst_en(x3503_sm_io_output_rst_en)
  );
  Counter_5 x3433 (
    .clock(x3433_clock),
    .reset(x3433_reset),
    .io_input_stops_0(x3433_io_input_stops_0),
    .io_input_reset(x3433_io_input_reset),
    .io_input_enable(x3433_io_input_enable),
    .io_output_counts_3(x3433_io_output_counts_3),
    .io_output_counts_2(x3433_io_output_counts_2),
    .io_output_counts_1(x3433_io_output_counts_1),
    .io_output_counts_0(x3433_io_output_counts_0),
    .io_output_done(x3433_io_output_done)
  );
  Innerpipe_10 x3466_sm (
    .clock(x3466_sm_clock),
    .reset(x3466_sm_reset),
    .io_input_enable(x3466_sm_io_input_enable),
    .io_input_ctr_done(x3466_sm_io_input_ctr_done),
    .io_input_rst(x3466_sm_io_input_rst),
    .io_output_done(x3466_sm_io_output_done),
    .io_output_ctr_inc(x3466_sm_io_output_ctr_inc),
    .io_output_rst_en(x3466_sm_io_output_rst_en)
  );
  Counter_5 x3469 (
    .clock(x3469_clock),
    .reset(x3469_reset),
    .io_input_stops_0(x3469_io_input_stops_0),
    .io_input_reset(x3469_io_input_reset),
    .io_input_enable(x3469_io_input_enable),
    .io_output_counts_3(x3469_io_output_counts_3),
    .io_output_counts_2(x3469_io_output_counts_2),
    .io_output_counts_1(x3469_io_output_counts_1),
    .io_output_counts_0(x3469_io_output_counts_0),
    .io_output_done(x3469_io_output_done)
  );
  Innerpipe_10 x3502_sm (
    .clock(x3502_sm_clock),
    .reset(x3502_sm_reset),
    .io_input_enable(x3502_sm_io_input_enable),
    .io_input_ctr_done(x3502_sm_io_input_ctr_done),
    .io_input_rst(x3502_sm_io_input_rst),
    .io_output_done(x3502_sm_io_output_done),
    .io_output_ctr_inc(x3502_sm_io_output_ctr_inc),
    .io_output_rst_en(x3502_sm_io_output_rst_en)
  );
  Innerpipe x3514_sm (
    .clock(x3514_sm_clock),
    .reset(x3514_sm_reset),
    .io_input_enable(x3514_sm_io_input_enable),
    .io_input_ctr_done(x3514_sm_io_input_ctr_done),
    .io_input_rst(x3514_sm_io_input_rst),
    .io_output_done(x3514_sm_io_output_done),
    .io_output_ctr_inc(x3514_sm_io_output_ctr_inc)
  );
  NBufFF_6 b1204_chain (
    .clock(b1204_chain_clock),
    .reset(b1204_chain_reset),
    .io_sEn_0(b1204_chain_io_sEn_0),
    .io_sEn_1(b1204_chain_io_sEn_1),
    .io_sEn_2(b1204_chain_io_sEn_2),
    .io_sEn_3(b1204_chain_io_sEn_3),
    .io_sEn_4(b1204_chain_io_sEn_4),
    .io_sDone_0(b1204_chain_io_sDone_0),
    .io_sDone_1(b1204_chain_io_sDone_1),
    .io_sDone_2(b1204_chain_io_sDone_2),
    .io_sDone_3(b1204_chain_io_sDone_3),
    .io_sDone_4(b1204_chain_io_sDone_4),
    .io_input_0_data(b1204_chain_io_input_0_data),
    .io_input_0_enable(b1204_chain_io_input_0_enable),
    .io_input_0_reset(b1204_chain_io_input_0_reset),
    .io_output_1_data(b1204_chain_io_output_1_data),
    .io_output_2_data(b1204_chain_io_output_2_data),
    .io_output_3_data(b1204_chain_io_output_3_data),
    .io_output_4_data(b1204_chain_io_output_4_data)
  );
  NBufFF_6 b1205_chain (
    .clock(b1205_chain_clock),
    .reset(b1205_chain_reset),
    .io_sEn_0(b1205_chain_io_sEn_0),
    .io_sEn_1(b1205_chain_io_sEn_1),
    .io_sEn_2(b1205_chain_io_sEn_2),
    .io_sEn_3(b1205_chain_io_sEn_3),
    .io_sEn_4(b1205_chain_io_sEn_4),
    .io_sDone_0(b1205_chain_io_sDone_0),
    .io_sDone_1(b1205_chain_io_sDone_1),
    .io_sDone_2(b1205_chain_io_sDone_2),
    .io_sDone_3(b1205_chain_io_sDone_3),
    .io_sDone_4(b1205_chain_io_sDone_4),
    .io_input_0_data(b1205_chain_io_input_0_data),
    .io_input_0_enable(b1205_chain_io_input_0_enable),
    .io_input_0_reset(b1205_chain_io_input_0_reset),
    .io_output_1_data(b1205_chain_io_output_1_data),
    .io_output_2_data(b1205_chain_io_output_2_data),
    .io_output_3_data(b1205_chain_io_output_3_data),
    .io_output_4_data(b1205_chain_io_output_4_data)
  );
  Innerpipe x3518_sm (
    .clock(x3518_sm_clock),
    .reset(x3518_sm_reset),
    .io_input_enable(x3518_sm_io_input_enable),
    .io_input_ctr_done(x3518_sm_io_input_ctr_done),
    .io_input_rst(x3518_sm_io_input_rst),
    .io_output_done(x3518_sm_io_output_done),
    .io_output_ctr_inc(x3518_sm_io_output_ctr_inc)
  );
  RetimeWrapper RetimeWrapper_1 (
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  SingleCounter_19 retime_counter (
    .clock(retime_counter_clock),
    .reset(retime_counter_reset),
    .io_input_reset(retime_counter_io_input_reset),
    .io_output_done(retime_counter_io_output_done)
  );
  RetimeWrapper RetimeWrapper_2 (
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 (
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 (
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 (
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 (
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 (
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper RetimeWrapper_8 (
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper RetimeWrapper_9 (
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper RetimeWrapper_10 (
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper RetimeWrapper_11 (
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper RetimeWrapper_12 (
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper RetimeWrapper_13 (
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper RetimeWrapper_14 (
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper RetimeWrapper_15 (
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper RetimeWrapper_16 (
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper RetimeWrapper_17 (
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper RetimeWrapper_18 (
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper RetimeWrapper_19 (
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper RetimeWrapper_20 (
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper RetimeWrapper_21 (
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper RetimeWrapper_22 (
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper RetimeWrapper_23 (
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper RetimeWrapper_24 (
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper RetimeWrapper_25 (
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper RetimeWrapper_26 (
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper RetimeWrapper_27 (
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper RetimeWrapper_28 (
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper RetimeWrapper_29 (
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper RetimeWrapper_30 (
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  SRFF done_latch (
    .clock(done_latch_clock),
    .reset(done_latch_reset),
    .io_input_set(done_latch_io_input_set),
    .io_input_reset(done_latch_io_input_reset),
    .io_input_asyn_reset(done_latch_io_input_asyn_reset),
    .io_output_data(done_latch_io_output_data)
  );
  RetimeWrapper RetimeWrapper_31 (
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper RetimeWrapper_32 (
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper RetimeWrapper_33 (
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper RetimeWrapper_34 (
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper RetimeWrapper_35 (
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper RetimeWrapper_36 (
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper RetimeWrapper_37 (
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper RetimeWrapper_38 (
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper RetimeWrapper_39 (
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper RetimeWrapper_40 (
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper RetimeWrapper_41 (
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper RetimeWrapper_42 (
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper RetimeWrapper_43 (
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper RetimeWrapper_44 (
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper RetimeWrapper_45 (
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper RetimeWrapper_46 (
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper RetimeWrapper_47 (
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper RetimeWrapper_48 (
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  RetimeWrapper RetimeWrapper_49 (
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper RetimeWrapper_50 (
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  RetimeWrapper RetimeWrapper_51 (
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  RetimeWrapper RetimeWrapper_52 (
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  RetimeWrapper RetimeWrapper_53 (
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  RetimeWrapper RetimeWrapper_54 (
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  RetimeWrapper RetimeWrapper_55 (
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  RetimeWrapper RetimeWrapper_56 (
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  RetimeWrapper RetimeWrapper_57 (
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  RetimeWrapper RetimeWrapper_58 (
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  RetimeWrapper RetimeWrapper_59 (
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper RetimeWrapper_60 (
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  RetimeWrapper RetimeWrapper_61 (
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  RetimeWrapper RetimeWrapper_62 (
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  RetimeWrapper RetimeWrapper_63 (
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  RetimeWrapper RetimeWrapper_64 (
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper RetimeWrapper_65 (
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  RetimeWrapper RetimeWrapper_66 (
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  RetimeWrapper RetimeWrapper_67 (
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  RetimeWrapper RetimeWrapper_68 (
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  RetimeWrapper RetimeWrapper_69 (
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  RetimeWrapper RetimeWrapper_70 (
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper RetimeWrapper_71 (
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  RetimeWrapper RetimeWrapper_72 (
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  RetimeWrapper RetimeWrapper_73 (
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  RetimeWrapper RetimeWrapper_74 (
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  RetimeWrapper RetimeWrapper_75 (
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  RetimeWrapper RetimeWrapper_76 (
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  RetimeWrapper RetimeWrapper_77 (
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  RetimeWrapper RetimeWrapper_78 (
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  RetimeWrapper RetimeWrapper_79 (
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  RetimeWrapper RetimeWrapper_80 (
    .clock(RetimeWrapper_80_clock),
    .reset(RetimeWrapper_80_reset),
    .io_flow(RetimeWrapper_80_io_flow),
    .io_in(RetimeWrapper_80_io_in),
    .io_out(RetimeWrapper_80_io_out)
  );
  RetimeWrapper RetimeWrapper_81 (
    .clock(RetimeWrapper_81_clock),
    .reset(RetimeWrapper_81_reset),
    .io_flow(RetimeWrapper_81_io_flow),
    .io_in(RetimeWrapper_81_io_in),
    .io_out(RetimeWrapper_81_io_out)
  );
  RetimeWrapper RetimeWrapper_82 (
    .clock(RetimeWrapper_82_clock),
    .reset(RetimeWrapper_82_reset),
    .io_flow(RetimeWrapper_82_io_flow),
    .io_in(RetimeWrapper_82_io_in),
    .io_out(RetimeWrapper_82_io_out)
  );
  RetimeWrapper RetimeWrapper_83 (
    .clock(RetimeWrapper_83_clock),
    .reset(RetimeWrapper_83_reset),
    .io_flow(RetimeWrapper_83_io_flow),
    .io_in(RetimeWrapper_83_io_in),
    .io_out(RetimeWrapper_83_io_out)
  );
  RetimeWrapper RetimeWrapper_84 (
    .clock(RetimeWrapper_84_clock),
    .reset(RetimeWrapper_84_reset),
    .io_flow(RetimeWrapper_84_io_flow),
    .io_in(RetimeWrapper_84_io_in),
    .io_out(RetimeWrapper_84_io_out)
  );
  RetimeWrapper RetimeWrapper_85 (
    .clock(RetimeWrapper_85_clock),
    .reset(RetimeWrapper_85_reset),
    .io_flow(RetimeWrapper_85_io_flow),
    .io_in(RetimeWrapper_85_io_in),
    .io_out(RetimeWrapper_85_io_out)
  );
  RetimeWrapper RetimeWrapper_86 (
    .clock(RetimeWrapper_86_clock),
    .reset(RetimeWrapper_86_reset),
    .io_flow(RetimeWrapper_86_io_flow),
    .io_in(RetimeWrapper_86_io_in),
    .io_out(RetimeWrapper_86_io_out)
  );
  RetimeWrapper RetimeWrapper_87 (
    .clock(RetimeWrapper_87_clock),
    .reset(RetimeWrapper_87_reset),
    .io_flow(RetimeWrapper_87_io_flow),
    .io_in(RetimeWrapper_87_io_in),
    .io_out(RetimeWrapper_87_io_out)
  );
  RetimeWrapper RetimeWrapper_88 (
    .clock(RetimeWrapper_88_clock),
    .reset(RetimeWrapper_88_reset),
    .io_flow(RetimeWrapper_88_io_flow),
    .io_in(RetimeWrapper_88_io_in),
    .io_out(RetimeWrapper_88_io_out)
  );
  RetimeWrapper RetimeWrapper_89 (
    .clock(RetimeWrapper_89_clock),
    .reset(RetimeWrapper_89_reset),
    .io_flow(RetimeWrapper_89_io_flow),
    .io_in(RetimeWrapper_89_io_in),
    .io_out(RetimeWrapper_89_io_out)
  );
  RetimeWrapper RetimeWrapper_90 (
    .clock(RetimeWrapper_90_clock),
    .reset(RetimeWrapper_90_reset),
    .io_flow(RetimeWrapper_90_io_flow),
    .io_in(RetimeWrapper_90_io_in),
    .io_out(RetimeWrapper_90_io_out)
  );
  RetimeWrapper RetimeWrapper_91 (
    .clock(RetimeWrapper_91_clock),
    .reset(RetimeWrapper_91_reset),
    .io_flow(RetimeWrapper_91_io_flow),
    .io_in(RetimeWrapper_91_io_in),
    .io_out(RetimeWrapper_91_io_out)
  );
  RetimeWrapper RetimeWrapper_92 (
    .clock(RetimeWrapper_92_clock),
    .reset(RetimeWrapper_92_reset),
    .io_flow(RetimeWrapper_92_io_flow),
    .io_in(RetimeWrapper_92_io_in),
    .io_out(RetimeWrapper_92_io_out)
  );
  RetimeWrapper RetimeWrapper_93 (
    .clock(RetimeWrapper_93_clock),
    .reset(RetimeWrapper_93_reset),
    .io_flow(RetimeWrapper_93_io_flow),
    .io_in(RetimeWrapper_93_io_in),
    .io_out(RetimeWrapper_93_io_out)
  );
  RetimeWrapper RetimeWrapper_94 (
    .clock(RetimeWrapper_94_clock),
    .reset(RetimeWrapper_94_reset),
    .io_flow(RetimeWrapper_94_io_flow),
    .io_in(RetimeWrapper_94_io_in),
    .io_out(RetimeWrapper_94_io_out)
  );
  RetimeWrapper RetimeWrapper_95 (
    .clock(RetimeWrapper_95_clock),
    .reset(RetimeWrapper_95_reset),
    .io_flow(RetimeWrapper_95_io_flow),
    .io_in(RetimeWrapper_95_io_in),
    .io_out(RetimeWrapper_95_io_out)
  );
  RetimeWrapper RetimeWrapper_96 (
    .clock(RetimeWrapper_96_clock),
    .reset(RetimeWrapper_96_reset),
    .io_flow(RetimeWrapper_96_io_flow),
    .io_in(RetimeWrapper_96_io_in),
    .io_out(RetimeWrapper_96_io_out)
  );
  RetimeWrapper RetimeWrapper_97 (
    .clock(RetimeWrapper_97_clock),
    .reset(RetimeWrapper_97_reset),
    .io_flow(RetimeWrapper_97_io_flow),
    .io_in(RetimeWrapper_97_io_in),
    .io_out(RetimeWrapper_97_io_out)
  );
  RetimeWrapper RetimeWrapper_98 (
    .clock(RetimeWrapper_98_clock),
    .reset(RetimeWrapper_98_reset),
    .io_flow(RetimeWrapper_98_io_flow),
    .io_in(RetimeWrapper_98_io_in),
    .io_out(RetimeWrapper_98_io_out)
  );
  RetimeWrapper RetimeWrapper_99 (
    .clock(RetimeWrapper_99_clock),
    .reset(RetimeWrapper_99_reset),
    .io_flow(RetimeWrapper_99_io_flow),
    .io_in(RetimeWrapper_99_io_in),
    .io_out(RetimeWrapper_99_io_out)
  );
  RetimeWrapper RetimeWrapper_100 (
    .clock(RetimeWrapper_100_clock),
    .reset(RetimeWrapper_100_reset),
    .io_flow(RetimeWrapper_100_io_flow),
    .io_in(RetimeWrapper_100_io_in),
    .io_out(RetimeWrapper_100_io_out)
  );
  RetimeWrapper RetimeWrapper_101 (
    .clock(RetimeWrapper_101_clock),
    .reset(RetimeWrapper_101_reset),
    .io_flow(RetimeWrapper_101_io_flow),
    .io_in(RetimeWrapper_101_io_in),
    .io_out(RetimeWrapper_101_io_out)
  );
  RetimeWrapper RetimeWrapper_102 (
    .clock(RetimeWrapper_102_clock),
    .reset(RetimeWrapper_102_reset),
    .io_flow(RetimeWrapper_102_io_flow),
    .io_in(RetimeWrapper_102_io_in),
    .io_out(RetimeWrapper_102_io_out)
  );
  RetimeWrapper RetimeWrapper_103 (
    .clock(RetimeWrapper_103_clock),
    .reset(RetimeWrapper_103_reset),
    .io_flow(RetimeWrapper_103_io_flow),
    .io_in(RetimeWrapper_103_io_in),
    .io_out(RetimeWrapper_103_io_out)
  );
  RetimeWrapper RetimeWrapper_104 (
    .clock(RetimeWrapper_104_clock),
    .reset(RetimeWrapper_104_reset),
    .io_flow(RetimeWrapper_104_io_flow),
    .io_in(RetimeWrapper_104_io_in),
    .io_out(RetimeWrapper_104_io_out)
  );
  RetimeWrapper RetimeWrapper_105 (
    .clock(RetimeWrapper_105_clock),
    .reset(RetimeWrapper_105_reset),
    .io_flow(RetimeWrapper_105_io_flow),
    .io_in(RetimeWrapper_105_io_in),
    .io_out(RetimeWrapper_105_io_out)
  );
  RetimeWrapper RetimeWrapper_106 (
    .clock(RetimeWrapper_106_clock),
    .reset(RetimeWrapper_106_reset),
    .io_flow(RetimeWrapper_106_io_flow),
    .io_in(RetimeWrapper_106_io_in),
    .io_out(RetimeWrapper_106_io_out)
  );
  RetimeWrapper RetimeWrapper_107 (
    .clock(RetimeWrapper_107_clock),
    .reset(RetimeWrapper_107_reset),
    .io_flow(RetimeWrapper_107_io_flow),
    .io_in(RetimeWrapper_107_io_in),
    .io_out(RetimeWrapper_107_io_out)
  );
  RetimeWrapper RetimeWrapper_108 (
    .clock(RetimeWrapper_108_clock),
    .reset(RetimeWrapper_108_reset),
    .io_flow(RetimeWrapper_108_io_flow),
    .io_in(RetimeWrapper_108_io_in),
    .io_out(RetimeWrapper_108_io_out)
  );
  RetimeWrapper RetimeWrapper_109 (
    .clock(RetimeWrapper_109_clock),
    .reset(RetimeWrapper_109_reset),
    .io_flow(RetimeWrapper_109_io_flow),
    .io_in(RetimeWrapper_109_io_in),
    .io_out(RetimeWrapper_109_io_out)
  );
  RetimeWrapper RetimeWrapper_110 (
    .clock(RetimeWrapper_110_clock),
    .reset(RetimeWrapper_110_reset),
    .io_flow(RetimeWrapper_110_io_flow),
    .io_in(RetimeWrapper_110_io_in),
    .io_out(RetimeWrapper_110_io_out)
  );
  RetimeWrapper RetimeWrapper_111 (
    .clock(RetimeWrapper_111_clock),
    .reset(RetimeWrapper_111_reset),
    .io_flow(RetimeWrapper_111_io_flow),
    .io_in(RetimeWrapper_111_io_in),
    .io_out(RetimeWrapper_111_io_out)
  );
  RetimeWrapper RetimeWrapper_112 (
    .clock(RetimeWrapper_112_clock),
    .reset(RetimeWrapper_112_reset),
    .io_flow(RetimeWrapper_112_io_flow),
    .io_in(RetimeWrapper_112_io_in),
    .io_out(RetimeWrapper_112_io_out)
  );
  RetimeWrapper RetimeWrapper_113 (
    .clock(RetimeWrapper_113_clock),
    .reset(RetimeWrapper_113_reset),
    .io_flow(RetimeWrapper_113_io_flow),
    .io_in(RetimeWrapper_113_io_in),
    .io_out(RetimeWrapper_113_io_out)
  );
  RetimeWrapper RetimeWrapper_114 (
    .clock(RetimeWrapper_114_clock),
    .reset(RetimeWrapper_114_reset),
    .io_flow(RetimeWrapper_114_io_flow),
    .io_in(RetimeWrapper_114_io_in),
    .io_out(RetimeWrapper_114_io_out)
  );
  RetimeWrapper RetimeWrapper_115 (
    .clock(RetimeWrapper_115_clock),
    .reset(RetimeWrapper_115_reset),
    .io_flow(RetimeWrapper_115_io_flow),
    .io_in(RetimeWrapper_115_io_in),
    .io_out(RetimeWrapper_115_io_out)
  );
  RetimeWrapper RetimeWrapper_116 (
    .clock(RetimeWrapper_116_clock),
    .reset(RetimeWrapper_116_reset),
    .io_flow(RetimeWrapper_116_io_flow),
    .io_in(RetimeWrapper_116_io_in),
    .io_out(RetimeWrapper_116_io_out)
  );
  RetimeWrapper RetimeWrapper_117 (
    .clock(RetimeWrapper_117_clock),
    .reset(RetimeWrapper_117_reset),
    .io_flow(RetimeWrapper_117_io_flow),
    .io_in(RetimeWrapper_117_io_in),
    .io_out(RetimeWrapper_117_io_out)
  );
  RetimeWrapper RetimeWrapper_118 (
    .clock(RetimeWrapper_118_clock),
    .reset(RetimeWrapper_118_reset),
    .io_flow(RetimeWrapper_118_io_flow),
    .io_in(RetimeWrapper_118_io_in),
    .io_out(RetimeWrapper_118_io_out)
  );
  RetimeWrapper RetimeWrapper_119 (
    .clock(RetimeWrapper_119_clock),
    .reset(RetimeWrapper_119_reset),
    .io_flow(RetimeWrapper_119_io_flow),
    .io_in(RetimeWrapper_119_io_in),
    .io_out(RetimeWrapper_119_io_out)
  );
  RetimeWrapper RetimeWrapper_120 (
    .clock(RetimeWrapper_120_clock),
    .reset(RetimeWrapper_120_reset),
    .io_flow(RetimeWrapper_120_io_flow),
    .io_in(RetimeWrapper_120_io_in),
    .io_out(RetimeWrapper_120_io_out)
  );
  RetimeWrapper RetimeWrapper_121 (
    .clock(RetimeWrapper_121_clock),
    .reset(RetimeWrapper_121_reset),
    .io_flow(RetimeWrapper_121_io_flow),
    .io_in(RetimeWrapper_121_io_in),
    .io_out(RetimeWrapper_121_io_out)
  );
  RetimeWrapper RetimeWrapper_122 (
    .clock(RetimeWrapper_122_clock),
    .reset(RetimeWrapper_122_reset),
    .io_flow(RetimeWrapper_122_io_flow),
    .io_in(RetimeWrapper_122_io_in),
    .io_out(RetimeWrapper_122_io_out)
  );
  RetimeWrapper RetimeWrapper_123 (
    .clock(RetimeWrapper_123_clock),
    .reset(RetimeWrapper_123_reset),
    .io_flow(RetimeWrapper_123_io_flow),
    .io_in(RetimeWrapper_123_io_in),
    .io_out(RetimeWrapper_123_io_out)
  );
  RetimeWrapper RetimeWrapper_124 (
    .clock(RetimeWrapper_124_clock),
    .reset(RetimeWrapper_124_reset),
    .io_flow(RetimeWrapper_124_io_flow),
    .io_in(RetimeWrapper_124_io_in),
    .io_out(RetimeWrapper_124_io_out)
  );
  RetimeWrapper RetimeWrapper_125 (
    .clock(RetimeWrapper_125_clock),
    .reset(RetimeWrapper_125_reset),
    .io_flow(RetimeWrapper_125_io_flow),
    .io_in(RetimeWrapper_125_io_in),
    .io_out(RetimeWrapper_125_io_out)
  );
  RetimeWrapper RetimeWrapper_126 (
    .clock(RetimeWrapper_126_clock),
    .reset(RetimeWrapper_126_reset),
    .io_flow(RetimeWrapper_126_io_flow),
    .io_in(RetimeWrapper_126_io_in),
    .io_out(RetimeWrapper_126_io_out)
  );
  RetimeWrapper RetimeWrapper_127 (
    .clock(RetimeWrapper_127_clock),
    .reset(RetimeWrapper_127_reset),
    .io_flow(RetimeWrapper_127_io_flow),
    .io_in(RetimeWrapper_127_io_in),
    .io_out(RetimeWrapper_127_io_out)
  );
  RetimeWrapper RetimeWrapper_128 (
    .clock(RetimeWrapper_128_clock),
    .reset(RetimeWrapper_128_reset),
    .io_flow(RetimeWrapper_128_io_flow),
    .io_in(RetimeWrapper_128_io_in),
    .io_out(RetimeWrapper_128_io_out)
  );
  RetimeWrapper RetimeWrapper_129 (
    .clock(RetimeWrapper_129_clock),
    .reset(RetimeWrapper_129_reset),
    .io_flow(RetimeWrapper_129_io_flow),
    .io_in(RetimeWrapper_129_io_in),
    .io_out(RetimeWrapper_129_io_out)
  );
  RetimeWrapper RetimeWrapper_130 (
    .clock(RetimeWrapper_130_clock),
    .reset(RetimeWrapper_130_reset),
    .io_flow(RetimeWrapper_130_io_flow),
    .io_in(RetimeWrapper_130_io_in),
    .io_out(RetimeWrapper_130_io_out)
  );
  RetimeWrapper RetimeWrapper_131 (
    .clock(RetimeWrapper_131_clock),
    .reset(RetimeWrapper_131_reset),
    .io_flow(RetimeWrapper_131_io_flow),
    .io_in(RetimeWrapper_131_io_in),
    .io_out(RetimeWrapper_131_io_out)
  );
  RetimeWrapper RetimeWrapper_132 (
    .clock(RetimeWrapper_132_clock),
    .reset(RetimeWrapper_132_reset),
    .io_flow(RetimeWrapper_132_io_flow),
    .io_in(RetimeWrapper_132_io_in),
    .io_out(RetimeWrapper_132_io_out)
  );
  RetimeWrapper RetimeWrapper_133 (
    .clock(RetimeWrapper_133_clock),
    .reset(RetimeWrapper_133_reset),
    .io_flow(RetimeWrapper_133_io_flow),
    .io_in(RetimeWrapper_133_io_in),
    .io_out(RetimeWrapper_133_io_out)
  );
  RetimeWrapper RetimeWrapper_134 (
    .clock(RetimeWrapper_134_clock),
    .reset(RetimeWrapper_134_reset),
    .io_flow(RetimeWrapper_134_io_flow),
    .io_in(RetimeWrapper_134_io_in),
    .io_out(RetimeWrapper_134_io_out)
  );
  RetimeWrapper RetimeWrapper_135 (
    .clock(RetimeWrapper_135_clock),
    .reset(RetimeWrapper_135_reset),
    .io_flow(RetimeWrapper_135_io_flow),
    .io_in(RetimeWrapper_135_io_in),
    .io_out(RetimeWrapper_135_io_out)
  );
  RetimeWrapper RetimeWrapper_136 (
    .clock(RetimeWrapper_136_clock),
    .reset(RetimeWrapper_136_reset),
    .io_flow(RetimeWrapper_136_io_flow),
    .io_in(RetimeWrapper_136_io_in),
    .io_out(RetimeWrapper_136_io_out)
  );
  RetimeWrapper RetimeWrapper_137 (
    .clock(RetimeWrapper_137_clock),
    .reset(RetimeWrapper_137_reset),
    .io_flow(RetimeWrapper_137_io_flow),
    .io_in(RetimeWrapper_137_io_in),
    .io_out(RetimeWrapper_137_io_out)
  );
  RetimeWrapper RetimeWrapper_138 (
    .clock(RetimeWrapper_138_clock),
    .reset(RetimeWrapper_138_reset),
    .io_flow(RetimeWrapper_138_io_flow),
    .io_in(RetimeWrapper_138_io_in),
    .io_out(RetimeWrapper_138_io_out)
  );
  RetimeWrapper RetimeWrapper_139 (
    .clock(RetimeWrapper_139_clock),
    .reset(RetimeWrapper_139_reset),
    .io_flow(RetimeWrapper_139_io_flow),
    .io_in(RetimeWrapper_139_io_in),
    .io_out(RetimeWrapper_139_io_out)
  );
  RetimeWrapper RetimeWrapper_140 (
    .clock(RetimeWrapper_140_clock),
    .reset(RetimeWrapper_140_reset),
    .io_flow(RetimeWrapper_140_io_flow),
    .io_in(RetimeWrapper_140_io_in),
    .io_out(RetimeWrapper_140_io_out)
  );
  RetimeWrapper RetimeWrapper_141 (
    .clock(RetimeWrapper_141_clock),
    .reset(RetimeWrapper_141_reset),
    .io_flow(RetimeWrapper_141_io_flow),
    .io_in(RetimeWrapper_141_io_in),
    .io_out(RetimeWrapper_141_io_out)
  );
  RetimeWrapper RetimeWrapper_142 (
    .clock(RetimeWrapper_142_clock),
    .reset(RetimeWrapper_142_reset),
    .io_flow(RetimeWrapper_142_io_flow),
    .io_in(RetimeWrapper_142_io_in),
    .io_out(RetimeWrapper_142_io_out)
  );
  RetimeWrapper RetimeWrapper_143 (
    .clock(RetimeWrapper_143_clock),
    .reset(RetimeWrapper_143_reset),
    .io_flow(RetimeWrapper_143_io_flow),
    .io_in(RetimeWrapper_143_io_in),
    .io_out(RetimeWrapper_143_io_out)
  );
  RetimeWrapper RetimeWrapper_144 (
    .clock(RetimeWrapper_144_clock),
    .reset(RetimeWrapper_144_reset),
    .io_flow(RetimeWrapper_144_io_flow),
    .io_in(RetimeWrapper_144_io_in),
    .io_out(RetimeWrapper_144_io_out)
  );
  RetimeWrapper RetimeWrapper_145 (
    .clock(RetimeWrapper_145_clock),
    .reset(RetimeWrapper_145_reset),
    .io_flow(RetimeWrapper_145_io_flow),
    .io_in(RetimeWrapper_145_io_in),
    .io_out(RetimeWrapper_145_io_out)
  );
  RetimeWrapper RetimeWrapper_146 (
    .clock(RetimeWrapper_146_clock),
    .reset(RetimeWrapper_146_reset),
    .io_flow(RetimeWrapper_146_io_flow),
    .io_in(RetimeWrapper_146_io_in),
    .io_out(RetimeWrapper_146_io_out)
  );
  RetimeWrapper RetimeWrapper_147 (
    .clock(RetimeWrapper_147_clock),
    .reset(RetimeWrapper_147_reset),
    .io_flow(RetimeWrapper_147_io_flow),
    .io_in(RetimeWrapper_147_io_in),
    .io_out(RetimeWrapper_147_io_out)
  );
  RetimeWrapper RetimeWrapper_148 (
    .clock(RetimeWrapper_148_clock),
    .reset(RetimeWrapper_148_reset),
    .io_flow(RetimeWrapper_148_io_flow),
    .io_in(RetimeWrapper_148_io_in),
    .io_out(RetimeWrapper_148_io_out)
  );
  RetimeWrapper RetimeWrapper_149 (
    .clock(RetimeWrapper_149_clock),
    .reset(RetimeWrapper_149_reset),
    .io_flow(RetimeWrapper_149_io_flow),
    .io_in(RetimeWrapper_149_io_in),
    .io_out(RetimeWrapper_149_io_out)
  );
  RetimeWrapper RetimeWrapper_150 (
    .clock(RetimeWrapper_150_clock),
    .reset(RetimeWrapper_150_reset),
    .io_flow(RetimeWrapper_150_io_flow),
    .io_in(RetimeWrapper_150_io_in),
    .io_out(RetimeWrapper_150_io_out)
  );
  RetimeWrapper RetimeWrapper_151 (
    .clock(RetimeWrapper_151_clock),
    .reset(RetimeWrapper_151_reset),
    .io_flow(RetimeWrapper_151_io_flow),
    .io_in(RetimeWrapper_151_io_in),
    .io_out(RetimeWrapper_151_io_out)
  );
  RetimeWrapper RetimeWrapper_152 (
    .clock(RetimeWrapper_152_clock),
    .reset(RetimeWrapper_152_reset),
    .io_flow(RetimeWrapper_152_io_flow),
    .io_in(RetimeWrapper_152_io_in),
    .io_out(RetimeWrapper_152_io_out)
  );
  RetimeWrapper RetimeWrapper_153 (
    .clock(RetimeWrapper_153_clock),
    .reset(RetimeWrapper_153_reset),
    .io_flow(RetimeWrapper_153_io_flow),
    .io_in(RetimeWrapper_153_io_in),
    .io_out(RetimeWrapper_153_io_out)
  );
  RetimeWrapper RetimeWrapper_154 (
    .clock(RetimeWrapper_154_clock),
    .reset(RetimeWrapper_154_reset),
    .io_flow(RetimeWrapper_154_io_flow),
    .io_in(RetimeWrapper_154_io_in),
    .io_out(RetimeWrapper_154_io_out)
  );
  RetimeWrapper RetimeWrapper_155 (
    .clock(RetimeWrapper_155_clock),
    .reset(RetimeWrapper_155_reset),
    .io_flow(RetimeWrapper_155_io_flow),
    .io_in(RetimeWrapper_155_io_in),
    .io_out(RetimeWrapper_155_io_out)
  );
  RetimeWrapper RetimeWrapper_156 (
    .clock(RetimeWrapper_156_clock),
    .reset(RetimeWrapper_156_reset),
    .io_flow(RetimeWrapper_156_io_flow),
    .io_in(RetimeWrapper_156_io_in),
    .io_out(RetimeWrapper_156_io_out)
  );
  RetimeWrapper RetimeWrapper_157 (
    .clock(RetimeWrapper_157_clock),
    .reset(RetimeWrapper_157_reset),
    .io_flow(RetimeWrapper_157_io_flow),
    .io_in(RetimeWrapper_157_io_in),
    .io_out(RetimeWrapper_157_io_out)
  );
  RetimeWrapper RetimeWrapper_158 (
    .clock(RetimeWrapper_158_clock),
    .reset(RetimeWrapper_158_reset),
    .io_flow(RetimeWrapper_158_io_flow),
    .io_in(RetimeWrapper_158_io_in),
    .io_out(RetimeWrapper_158_io_out)
  );
  RetimeWrapper RetimeWrapper_159 (
    .clock(RetimeWrapper_159_clock),
    .reset(RetimeWrapper_159_reset),
    .io_flow(RetimeWrapper_159_io_flow),
    .io_in(RetimeWrapper_159_io_in),
    .io_out(RetimeWrapper_159_io_out)
  );
  RetimeWrapper RetimeWrapper_160 (
    .clock(RetimeWrapper_160_clock),
    .reset(RetimeWrapper_160_reset),
    .io_flow(RetimeWrapper_160_io_flow),
    .io_in(RetimeWrapper_160_io_in),
    .io_out(RetimeWrapper_160_io_out)
  );
  RetimeWrapper RetimeWrapper_161 (
    .clock(RetimeWrapper_161_clock),
    .reset(RetimeWrapper_161_reset),
    .io_flow(RetimeWrapper_161_io_flow),
    .io_in(RetimeWrapper_161_io_in),
    .io_out(RetimeWrapper_161_io_out)
  );
  RetimeWrapper RetimeWrapper_162 (
    .clock(RetimeWrapper_162_clock),
    .reset(RetimeWrapper_162_reset),
    .io_flow(RetimeWrapper_162_io_flow),
    .io_in(RetimeWrapper_162_io_in),
    .io_out(RetimeWrapper_162_io_out)
  );
  RetimeWrapper RetimeWrapper_163 (
    .clock(RetimeWrapper_163_clock),
    .reset(RetimeWrapper_163_reset),
    .io_flow(RetimeWrapper_163_io_flow),
    .io_in(RetimeWrapper_163_io_in),
    .io_out(RetimeWrapper_163_io_out)
  );
  RetimeWrapper RetimeWrapper_164 (
    .clock(RetimeWrapper_164_clock),
    .reset(RetimeWrapper_164_reset),
    .io_flow(RetimeWrapper_164_io_flow),
    .io_in(RetimeWrapper_164_io_in),
    .io_out(RetimeWrapper_164_io_out)
  );
  RetimeWrapper RetimeWrapper_165 (
    .clock(RetimeWrapper_165_clock),
    .reset(RetimeWrapper_165_reset),
    .io_flow(RetimeWrapper_165_io_flow),
    .io_in(RetimeWrapper_165_io_in),
    .io_out(RetimeWrapper_165_io_out)
  );
  RetimeWrapper RetimeWrapper_166 (
    .clock(RetimeWrapper_166_clock),
    .reset(RetimeWrapper_166_reset),
    .io_flow(RetimeWrapper_166_io_flow),
    .io_in(RetimeWrapper_166_io_in),
    .io_out(RetimeWrapper_166_io_out)
  );
  RetimeWrapper RetimeWrapper_167 (
    .clock(RetimeWrapper_167_clock),
    .reset(RetimeWrapper_167_reset),
    .io_flow(RetimeWrapper_167_io_flow),
    .io_in(RetimeWrapper_167_io_in),
    .io_out(RetimeWrapper_167_io_out)
  );
  RetimeWrapper RetimeWrapper_168 (
    .clock(RetimeWrapper_168_clock),
    .reset(RetimeWrapper_168_reset),
    .io_flow(RetimeWrapper_168_io_flow),
    .io_in(RetimeWrapper_168_io_in),
    .io_out(RetimeWrapper_168_io_out)
  );
  RetimeWrapper RetimeWrapper_169 (
    .clock(RetimeWrapper_169_clock),
    .reset(RetimeWrapper_169_reset),
    .io_flow(RetimeWrapper_169_io_flow),
    .io_in(RetimeWrapper_169_io_in),
    .io_out(RetimeWrapper_169_io_out)
  );
  RetimeWrapper RetimeWrapper_170 (
    .clock(RetimeWrapper_170_clock),
    .reset(RetimeWrapper_170_reset),
    .io_flow(RetimeWrapper_170_io_flow),
    .io_in(RetimeWrapper_170_io_in),
    .io_out(RetimeWrapper_170_io_out)
  );
  RetimeWrapper RetimeWrapper_171 (
    .clock(RetimeWrapper_171_clock),
    .reset(RetimeWrapper_171_reset),
    .io_flow(RetimeWrapper_171_io_flow),
    .io_in(RetimeWrapper_171_io_in),
    .io_out(RetimeWrapper_171_io_out)
  );
  RetimeWrapper RetimeWrapper_172 (
    .clock(RetimeWrapper_172_clock),
    .reset(RetimeWrapper_172_reset),
    .io_flow(RetimeWrapper_172_io_flow),
    .io_in(RetimeWrapper_172_io_in),
    .io_out(RetimeWrapper_172_io_out)
  );
  RetimeWrapper RetimeWrapper_173 (
    .clock(RetimeWrapper_173_clock),
    .reset(RetimeWrapper_173_reset),
    .io_flow(RetimeWrapper_173_io_flow),
    .io_in(RetimeWrapper_173_io_in),
    .io_out(RetimeWrapper_173_io_out)
  );
  RetimeWrapper RetimeWrapper_174 (
    .clock(RetimeWrapper_174_clock),
    .reset(RetimeWrapper_174_reset),
    .io_flow(RetimeWrapper_174_io_flow),
    .io_in(RetimeWrapper_174_io_in),
    .io_out(RetimeWrapper_174_io_out)
  );
  RetimeWrapper RetimeWrapper_175 (
    .clock(RetimeWrapper_175_clock),
    .reset(RetimeWrapper_175_reset),
    .io_flow(RetimeWrapper_175_io_flow),
    .io_in(RetimeWrapper_175_io_in),
    .io_out(RetimeWrapper_175_io_out)
  );
  RetimeWrapper RetimeWrapper_176 (
    .clock(RetimeWrapper_176_clock),
    .reset(RetimeWrapper_176_reset),
    .io_flow(RetimeWrapper_176_io_flow),
    .io_in(RetimeWrapper_176_io_in),
    .io_out(RetimeWrapper_176_io_out)
  );
  RetimeWrapper RetimeWrapper_177 (
    .clock(RetimeWrapper_177_clock),
    .reset(RetimeWrapper_177_reset),
    .io_flow(RetimeWrapper_177_io_flow),
    .io_in(RetimeWrapper_177_io_in),
    .io_out(RetimeWrapper_177_io_out)
  );
  RetimeWrapper RetimeWrapper_178 (
    .clock(RetimeWrapper_178_clock),
    .reset(RetimeWrapper_178_reset),
    .io_flow(RetimeWrapper_178_io_flow),
    .io_in(RetimeWrapper_178_io_in),
    .io_out(RetimeWrapper_178_io_out)
  );
  RetimeWrapper RetimeWrapper_179 (
    .clock(RetimeWrapper_179_clock),
    .reset(RetimeWrapper_179_reset),
    .io_flow(RetimeWrapper_179_io_flow),
    .io_in(RetimeWrapper_179_io_in),
    .io_out(RetimeWrapper_179_io_out)
  );
  RetimeWrapper RetimeWrapper_180 (
    .clock(RetimeWrapper_180_clock),
    .reset(RetimeWrapper_180_reset),
    .io_flow(RetimeWrapper_180_io_flow),
    .io_in(RetimeWrapper_180_io_in),
    .io_out(RetimeWrapper_180_io_out)
  );
  RetimeWrapper RetimeWrapper_181 (
    .clock(RetimeWrapper_181_clock),
    .reset(RetimeWrapper_181_reset),
    .io_flow(RetimeWrapper_181_io_flow),
    .io_in(RetimeWrapper_181_io_in),
    .io_out(RetimeWrapper_181_io_out)
  );
  RetimeWrapper RetimeWrapper_182 (
    .clock(RetimeWrapper_182_clock),
    .reset(RetimeWrapper_182_reset),
    .io_flow(RetimeWrapper_182_io_flow),
    .io_in(RetimeWrapper_182_io_in),
    .io_out(RetimeWrapper_182_io_out)
  );
  RetimeWrapper RetimeWrapper_183 (
    .clock(RetimeWrapper_183_clock),
    .reset(RetimeWrapper_183_reset),
    .io_flow(RetimeWrapper_183_io_flow),
    .io_in(RetimeWrapper_183_io_in),
    .io_out(RetimeWrapper_183_io_out)
  );
  RetimeWrapper RetimeWrapper_184 (
    .clock(RetimeWrapper_184_clock),
    .reset(RetimeWrapper_184_reset),
    .io_flow(RetimeWrapper_184_io_flow),
    .io_in(RetimeWrapper_184_io_in),
    .io_out(RetimeWrapper_184_io_out)
  );
  RetimeWrapper RetimeWrapper_185 (
    .clock(RetimeWrapper_185_clock),
    .reset(RetimeWrapper_185_reset),
    .io_flow(RetimeWrapper_185_io_flow),
    .io_in(RetimeWrapper_185_io_in),
    .io_out(RetimeWrapper_185_io_out)
  );
  RetimeWrapper RetimeWrapper_186 (
    .clock(RetimeWrapper_186_clock),
    .reset(RetimeWrapper_186_reset),
    .io_flow(RetimeWrapper_186_io_flow),
    .io_in(RetimeWrapper_186_io_in),
    .io_out(RetimeWrapper_186_io_out)
  );
  RetimeWrapper RetimeWrapper_187 (
    .clock(RetimeWrapper_187_clock),
    .reset(RetimeWrapper_187_reset),
    .io_flow(RetimeWrapper_187_io_flow),
    .io_in(RetimeWrapper_187_io_in),
    .io_out(RetimeWrapper_187_io_out)
  );
  RetimeWrapper RetimeWrapper_188 (
    .clock(RetimeWrapper_188_clock),
    .reset(RetimeWrapper_188_reset),
    .io_flow(RetimeWrapper_188_io_flow),
    .io_in(RetimeWrapper_188_io_in),
    .io_out(RetimeWrapper_188_io_out)
  );
  RetimeWrapper RetimeWrapper_189 (
    .clock(RetimeWrapper_189_clock),
    .reset(RetimeWrapper_189_reset),
    .io_flow(RetimeWrapper_189_io_flow),
    .io_in(RetimeWrapper_189_io_in),
    .io_out(RetimeWrapper_189_io_out)
  );
  RetimeWrapper RetimeWrapper_190 (
    .clock(RetimeWrapper_190_clock),
    .reset(RetimeWrapper_190_reset),
    .io_flow(RetimeWrapper_190_io_flow),
    .io_in(RetimeWrapper_190_io_in),
    .io_out(RetimeWrapper_190_io_out)
  );
  RetimeWrapper RetimeWrapper_191 (
    .clock(RetimeWrapper_191_clock),
    .reset(RetimeWrapper_191_reset),
    .io_flow(RetimeWrapper_191_io_flow),
    .io_in(RetimeWrapper_191_io_in),
    .io_out(RetimeWrapper_191_io_out)
  );
  RetimeWrapper RetimeWrapper_192 (
    .clock(RetimeWrapper_192_clock),
    .reset(RetimeWrapper_192_reset),
    .io_flow(RetimeWrapper_192_io_flow),
    .io_in(RetimeWrapper_192_io_in),
    .io_out(RetimeWrapper_192_io_out)
  );
  RetimeWrapper RetimeWrapper_193 (
    .clock(RetimeWrapper_193_clock),
    .reset(RetimeWrapper_193_reset),
    .io_flow(RetimeWrapper_193_io_flow),
    .io_in(RetimeWrapper_193_io_in),
    .io_out(RetimeWrapper_193_io_out)
  );
  RetimeWrapper RetimeWrapper_194 (
    .clock(RetimeWrapper_194_clock),
    .reset(RetimeWrapper_194_reset),
    .io_flow(RetimeWrapper_194_io_flow),
    .io_in(RetimeWrapper_194_io_in),
    .io_out(RetimeWrapper_194_io_out)
  );
  RetimeWrapper RetimeWrapper_195 (
    .clock(RetimeWrapper_195_clock),
    .reset(RetimeWrapper_195_reset),
    .io_flow(RetimeWrapper_195_io_flow),
    .io_in(RetimeWrapper_195_io_in),
    .io_out(RetimeWrapper_195_io_out)
  );
  RetimeWrapper RetimeWrapper_196 (
    .clock(RetimeWrapper_196_clock),
    .reset(RetimeWrapper_196_reset),
    .io_flow(RetimeWrapper_196_io_flow),
    .io_in(RetimeWrapper_196_io_in),
    .io_out(RetimeWrapper_196_io_out)
  );
  RetimeWrapper RetimeWrapper_197 (
    .clock(RetimeWrapper_197_clock),
    .reset(RetimeWrapper_197_reset),
    .io_flow(RetimeWrapper_197_io_flow),
    .io_in(RetimeWrapper_197_io_in),
    .io_out(RetimeWrapper_197_io_out)
  );
  RetimeWrapper RetimeWrapper_198 (
    .clock(RetimeWrapper_198_clock),
    .reset(RetimeWrapper_198_reset),
    .io_flow(RetimeWrapper_198_io_flow),
    .io_in(RetimeWrapper_198_io_in),
    .io_out(RetimeWrapper_198_io_out)
  );
  RetimeWrapper RetimeWrapper_199 (
    .clock(RetimeWrapper_199_clock),
    .reset(RetimeWrapper_199_reset),
    .io_flow(RetimeWrapper_199_io_flow),
    .io_in(RetimeWrapper_199_io_in),
    .io_out(RetimeWrapper_199_io_out)
  );
  RetimeWrapper RetimeWrapper_200 (
    .clock(RetimeWrapper_200_clock),
    .reset(RetimeWrapper_200_reset),
    .io_flow(RetimeWrapper_200_io_flow),
    .io_in(RetimeWrapper_200_io_in),
    .io_out(RetimeWrapper_200_io_out)
  );
  RetimeWrapper RetimeWrapper_201 (
    .clock(RetimeWrapper_201_clock),
    .reset(RetimeWrapper_201_reset),
    .io_flow(RetimeWrapper_201_io_flow),
    .io_in(RetimeWrapper_201_io_in),
    .io_out(RetimeWrapper_201_io_out)
  );
  RetimeWrapper RetimeWrapper_202 (
    .clock(RetimeWrapper_202_clock),
    .reset(RetimeWrapper_202_reset),
    .io_flow(RetimeWrapper_202_io_flow),
    .io_in(RetimeWrapper_202_io_in),
    .io_out(RetimeWrapper_202_io_out)
  );
  RetimeWrapper RetimeWrapper_203 (
    .clock(RetimeWrapper_203_clock),
    .reset(RetimeWrapper_203_reset),
    .io_flow(RetimeWrapper_203_io_flow),
    .io_in(RetimeWrapper_203_io_in),
    .io_out(RetimeWrapper_203_io_out)
  );
  RetimeWrapper RetimeWrapper_204 (
    .clock(RetimeWrapper_204_clock),
    .reset(RetimeWrapper_204_reset),
    .io_flow(RetimeWrapper_204_io_flow),
    .io_in(RetimeWrapper_204_io_in),
    .io_out(RetimeWrapper_204_io_out)
  );
  RetimeWrapper RetimeWrapper_205 (
    .clock(RetimeWrapper_205_clock),
    .reset(RetimeWrapper_205_reset),
    .io_flow(RetimeWrapper_205_io_flow),
    .io_in(RetimeWrapper_205_io_in),
    .io_out(RetimeWrapper_205_io_out)
  );
  RetimeWrapper RetimeWrapper_206 (
    .clock(RetimeWrapper_206_clock),
    .reset(RetimeWrapper_206_reset),
    .io_flow(RetimeWrapper_206_io_flow),
    .io_in(RetimeWrapper_206_io_in),
    .io_out(RetimeWrapper_206_io_out)
  );
  RetimeWrapper RetimeWrapper_207 (
    .clock(RetimeWrapper_207_clock),
    .reset(RetimeWrapper_207_reset),
    .io_flow(RetimeWrapper_207_io_flow),
    .io_in(RetimeWrapper_207_io_in),
    .io_out(RetimeWrapper_207_io_out)
  );
  RetimeWrapper RetimeWrapper_208 (
    .clock(RetimeWrapper_208_clock),
    .reset(RetimeWrapper_208_reset),
    .io_flow(RetimeWrapper_208_io_flow),
    .io_in(RetimeWrapper_208_io_in),
    .io_out(RetimeWrapper_208_io_out)
  );
  RetimeWrapper RetimeWrapper_209 (
    .clock(RetimeWrapper_209_clock),
    .reset(RetimeWrapper_209_reset),
    .io_flow(RetimeWrapper_209_io_flow),
    .io_in(RetimeWrapper_209_io_in),
    .io_out(RetimeWrapper_209_io_out)
  );
  RetimeWrapper RetimeWrapper_210 (
    .clock(RetimeWrapper_210_clock),
    .reset(RetimeWrapper_210_reset),
    .io_flow(RetimeWrapper_210_io_flow),
    .io_in(RetimeWrapper_210_io_in),
    .io_out(RetimeWrapper_210_io_out)
  );
  RetimeWrapper RetimeWrapper_211 (
    .clock(RetimeWrapper_211_clock),
    .reset(RetimeWrapper_211_reset),
    .io_flow(RetimeWrapper_211_io_flow),
    .io_in(RetimeWrapper_211_io_in),
    .io_out(RetimeWrapper_211_io_out)
  );
  RetimeWrapper RetimeWrapper_212 (
    .clock(RetimeWrapper_212_clock),
    .reset(RetimeWrapper_212_reset),
    .io_flow(RetimeWrapper_212_io_flow),
    .io_in(RetimeWrapper_212_io_in),
    .io_out(RetimeWrapper_212_io_out)
  );
  assign _T_1601 = x3175_valid_stops_0 | reset;
  assign _T_1610 = x3238_valid_stops_0 | reset;
  assign _T_1619 = x3302_valid_stops_0 | reset;
  assign _T_1628 = x3365_valid_stops_0 | reset;
  assign _T_1660 = b1204_chain_io_output_1_data;
  assign _T_1662 = b1204_chain_io_output_2_data;
  assign _T_1664 = b1204_chain_io_output_3_data;
  assign _T_1668 = b1205_chain_io_output_1_data;
  assign _T_1670 = b1205_chain_io_output_2_data;
  assign _T_1672 = b1205_chain_io_output_3_data;
  assign _T_1674 = b1205_chain_io_output_4_data;
  assign _T_1675 = RootController_en & retime_released;
  assign _T_1678 = retime_released ? RootController_sm_io_output_done : 1'h0;
  assign _T_1679 = ~ _T_1678;
  assign _T_1688 = _T_1678 & _T_1682;
  assign _T_1697 = io_done == 1'h0;
  assign _T_1698 = io_enable & _T_1697;
  assign _T_1711 = $signed(x3153_number);
  assign _T_1737 = x3153_number[31];
  assign _T_1739 = {_T_1737,x3153_number};
  assign _T_1753 = _T_1724_number - 33'h0;
  assign _T_1754 = $unsigned(_T_1753);
  assign _T_1755 = _T_1754[32:0];
  assign _T_1774 = _T_1722_number[31:0];
  assign _T_1780 = $signed(x35150_range_number);
  assign _T_1782 = $signed(_T_1780) / $signed(32'sh80);
  assign _T_1784 = $unsigned(_T_1782);
  assign _GEN_8 = x35150_range_number % 32'h80;
  assign _T_1806 = _GEN_8[31:0];
  assign _T_1881 = _T_1805_number[31:0];
  assign x35150_evenfit = x35150_leftover_number == 32'h0;
  assign x35150_adjustment = x35150_evenfit ? 1'h0 : 1'h1;
  assign _T_1928 = {31'h0,_T_1911_number};
  assign _T_1947 = {1'h0,x35150_hops_number};
  assign _T_1960 = {1'h0,_T_1909_number};
  assign _T_1961 = _T_1932_number + _T_1934_number;
  assign _T_1962 = _T_1961[32:0];
  assign _T_1976 = _T_1930_number[31:0];
  assign _T_1978 = x3515_en & retime_released;
  assign _T_1981 = retime_released ? x3515_sm_io_output_done : 1'h0;
  assign _T_1982 = ~ _T_1981;
  assign _T_1991 = _T_1981 & _T_1985;
  assign _T_1992 = ~ x3515_done;
  assign _T_1996 = x3515_sm_io_output_ctr_inc;
  assign _T_1999 = retime_released ? x3515_rst_en : 1'h0;
  assign _T_2100 = $signed(_T_2075_number);
  assign _T_2101 = $signed(_T_2077_number);
  assign _T_2102 = $signed(_T_2100) < $signed(_T_2101);
  assign _T_2237 = $signed(_T_2212_number);
  assign _T_2238 = $signed(_T_2214_number);
  assign _T_2239 = $signed(_T_2237) < $signed(_T_2238);
  assign _T_2282 = retime_released ? _T_2280 : 1'h0;
  assign _T_2283 = ~ x3174_done;
  assign _T_2289 = retime_released ? _T_2287 : 1'h0;
  assign _T_2290 = _T_2282 & _T_2289;
  assign _T_2296 = retime_released ? _T_2294 : 1'h0;
  assign _T_2302 = retime_released ? _T_2300 : 1'h0;
  assign _T_2303 = ~ x3301_done;
  assign _T_2309 = retime_released ? _T_2307 : 1'h0;
  assign _T_2310 = _T_2302 & _T_2309;
  assign _T_2316 = retime_released ? _T_2314 : 1'h0;
  assign _T_2322 = retime_released ? _T_2320 : 1'h0;
  assign _T_2323 = ~ x3428_done;
  assign _T_2329 = retime_released ? _T_2327 : 1'h0;
  assign _T_2330 = _T_2322 & _T_2329;
  assign _T_2336 = retime_released ? _T_2334 : 1'h0;
  assign _T_2342 = retime_released ? _T_2340 : 1'h0;
  assign _T_2343 = ~ x3503_done;
  assign _T_2349 = retime_released ? _T_2347 : 1'h0;
  assign _T_2350 = _T_2342 & _T_2349;
  assign _T_2356 = retime_released ? _T_2354 : 1'h0;
  assign _T_2362 = retime_released ? _T_2360 : 1'h0;
  assign _T_2363 = ~ x3514_done;
  assign _T_2369 = retime_released ? _T_2367 : 1'h0;
  assign _T_2370 = _T_2362 & _T_2369;
  assign _T_2376 = retime_released ? _T_2374 : 1'h0;
  assign _T_2396 = retime_released ? _T_2394 : 1'h0;
  assign _T_2423 = _T_2398_number == 32'h0;
  assign _T_2424 = _T_2396 | _T_2423;
  assign _T_2426 = x3518_en & retime_released;
  assign _T_2429 = retime_released ? x3518_sm_io_output_done : 1'h0;
  assign _T_2430 = ~ _T_2429;
  assign _T_2439 = _T_2429 & _T_2433;
  assign _T_2441 = ~ x3518_done;
  assign _T_2442 = x3518_sm_io_output_ctr_inc & _T_2441;
  assign _T_2443 = ~ x3518_ctr_trivial;
  assign _T_2444 = _T_2442 & _T_2443;
  assign _T_2445 = ~ x3518_sm_io_output_ctr_inc;
  assign _T_2454 = x3518_sm_io_output_ctr_inc & _T_2448;
  assign _T_2460 = retime_released ? _T_2458 : 1'h0;
  assign _T_2468 = retime_released ? _T_2466 : 1'h0;
  assign _T_2478 = retime_released ? _T_2476 : 1'h0;
  assign _T_2485 = retime_released ? _T_2483 : 1'h0;
  assign _T_2486 = _T_2478 & _T_2485;
  assign _T_2492 = retime_released ? _T_2490 : 1'h0;
  assign _T_2498 = retime_released ? _T_2496 : 1'h0;
  assign _T_2505 = retime_released ? _T_2503 : 1'h0;
  assign _T_2506 = _T_2498 & _T_2505;
  assign _T_2512 = retime_released ? _T_2510 : 1'h0;
  assign _T_2513 = $unsigned(x3154_0);
  assign _T_2514 = $unsigned(x3154_1);
  assign _T_2517 = x3174_en & retime_released;
  assign _T_2520 = retime_released ? x3174_sm_io_output_done : 1'h0;
  assign _T_2521 = ~ _T_2520;
  assign _T_2530 = _T_2520 & _T_2524;
  assign _T_2543 = retime_released ? _T_2541 : 1'h0;
  assign _T_2551 = retime_released ? _T_2549 : 1'h0;
  assign _T_2552 = ~ x3167_done;
  assign _T_2558 = retime_released ? _T_2556 : 1'h0;
  assign _T_2559 = _T_2551 & _T_2558;
  assign _T_2565 = retime_released ? _T_2563 : 1'h0;
  assign _T_2571 = retime_released ? _T_2569 : 1'h0;
  assign _T_2572 = ~ x3173_done;
  assign _T_2578 = retime_released ? _T_2576 : 1'h0;
  assign _T_2579 = _T_2571 & _T_2578;
  assign _T_2585 = retime_released ? _T_2583 : 1'h0;
  assign _T_2587 = x3301_en & retime_released;
  assign _T_2590 = retime_released ? x3301_sm_io_output_done : 1'h0;
  assign _T_2591 = ~ _T_2590;
  assign _T_2600 = _T_2590 & _T_2594;
  assign _T_2613 = retime_released ? _T_2611 : 1'h0;
  assign _T_2621 = retime_released ? _T_2619 : 1'h0;
  assign _T_2622 = ~ x3237_done;
  assign _T_2628 = retime_released ? _T_2626 : 1'h0;
  assign _T_2629 = _T_2621 & _T_2628;
  assign _T_2635 = retime_released ? _T_2633 : 1'h0;
  assign _T_2641 = retime_released ? _T_2639 : 1'h0;
  assign _T_2642 = ~ x3300_done;
  assign _T_2648 = retime_released ? _T_2646 : 1'h0;
  assign _T_2649 = _T_2641 & _T_2648;
  assign _T_2655 = retime_released ? _T_2653 : 1'h0;
  assign _T_2657 = x3428_en & retime_released;
  assign _T_2660 = retime_released ? x3428_sm_io_output_done : 1'h0;
  assign _T_2661 = ~ _T_2660;
  assign _T_2670 = _T_2660 & _T_2664;
  assign _T_2683 = retime_released ? _T_2681 : 1'h0;
  assign _T_2691 = retime_released ? _T_2689 : 1'h0;
  assign _T_2692 = ~ x3364_done;
  assign _T_2698 = retime_released ? _T_2696 : 1'h0;
  assign _T_2699 = _T_2691 & _T_2698;
  assign _T_2705 = retime_released ? _T_2703 : 1'h0;
  assign _T_2711 = retime_released ? _T_2709 : 1'h0;
  assign _T_2712 = ~ x3427_done;
  assign _T_2718 = retime_released ? _T_2716 : 1'h0;
  assign _T_2719 = _T_2711 & _T_2718;
  assign _T_2725 = retime_released ? _T_2723 : 1'h0;
  assign _T_2729 = x3503_en & retime_released;
  assign _T_2732 = retime_released ? x3503_sm_io_output_done : 1'h0;
  assign _T_2733 = ~ _T_2732;
  assign _T_2742 = _T_2732 & _T_2736;
  assign _T_2755 = retime_released ? _T_2753 : 1'h0;
  assign _T_2763 = retime_released ? _T_2761 : 1'h0;
  assign _T_2764 = ~ x3466_done;
  assign _T_2770 = retime_released ? _T_2768 : 1'h0;
  assign _T_2771 = _T_2763 & _T_2770;
  assign _T_2777 = retime_released ? _T_2775 : 1'h0;
  assign _T_2783 = retime_released ? _T_2781 : 1'h0;
  assign _T_2784 = ~ x3502_done;
  assign _T_2790 = retime_released ? _T_2788 : 1'h0;
  assign _T_2791 = _T_2783 & _T_2790;
  assign _T_2797 = retime_released ? _T_2795 : 1'h0;
  assign _T_2799 = x3514_en & retime_released;
  assign _T_2802 = retime_released ? x3514_sm_io_output_done : 1'h0;
  assign _T_2803 = ~ _T_2802;
  assign _T_2812 = _T_2802 & _T_2806;
  assign _T_2818 = ~ x3514_sm_io_output_ctr_inc;
  assign _T_2827 = x3514_sm_io_output_ctr_inc & _T_2821;
  assign _T_2833 = retime_released ? _T_2831 : 1'h0;
  assign _T_2846 = x3237_en & retime_released;
  assign _T_2848 = x3237_sm_io_output_done;
  assign _T_2861 = retime_released ? _T_2859 : 1'h0;
  assign _T_2869 = retime_released ? _T_2867 : 1'h0;
  assign _T_2870 = ~ x3208_done;
  assign _T_2876 = retime_released ? _T_2874 : 1'h0;
  assign _T_2877 = _T_2869 & _T_2876;
  assign _T_2878 = x3208_base_en & x3175_ready;
  assign _T_2879 = ~ x3176_io_full;
  assign _T_2885 = retime_released ? _T_2883 : 1'h0;
  assign _T_2886 = ~ b1204_chain_read_1;
  assign _T_2887 = _T_2885 | _T_2886;
  assign _T_2888 = _T_2878 & _T_2887;
  assign _T_2894 = retime_released ? _T_2892 : 1'h0;
  assign _T_2900 = retime_released ? _T_2898 : 1'h0;
  assign _T_2901 = ~ x3236_done;
  assign _T_2907 = retime_released ? _T_2905 : 1'h0;
  assign _T_2908 = _T_2900 & _T_2907;
  assign _T_2914 = retime_released ? _T_2912 : 1'h0;
  assign _T_2915 = x3300_en & retime_released;
  assign _T_2917 = x3300_sm_io_output_done;
  assign _T_2930 = retime_released ? _T_2928 : 1'h0;
  assign _T_2938 = retime_released ? _T_2936 : 1'h0;
  assign _T_2939 = ~ x3271_done;
  assign _T_2945 = retime_released ? _T_2943 : 1'h0;
  assign _T_2946 = _T_2938 & _T_2945;
  assign _T_2947 = x3271_base_en & x3238_ready;
  assign _T_2948 = ~ x3239_io_full;
  assign _T_2954 = retime_released ? _T_2952 : 1'h0;
  assign _T_2955 = ~ b1205_chain_read_1;
  assign _T_2956 = _T_2954 | _T_2955;
  assign _T_2957 = _T_2947 & _T_2956;
  assign _T_2963 = retime_released ? _T_2961 : 1'h0;
  assign _T_2969 = retime_released ? _T_2967 : 1'h0;
  assign _T_2970 = ~ x3299_done;
  assign _T_2976 = retime_released ? _T_2974 : 1'h0;
  assign _T_2977 = _T_2969 & _T_2976;
  assign _T_2983 = retime_released ? _T_2981 : 1'h0;
  assign _T_2984 = x3208_en & retime_released;
  assign _T_2986 = x3175_ready & _T_2879;
  assign _T_2987 = x3208_sm_io_output_done & _T_2986;
  assign _T_2990 = x3208_sm_io_output_ctr_inc & _T_2870;
  assign _T_2991 = ~ x3208_ctr_trivial;
  assign _T_2992 = _T_2990 & _T_2991;
  assign _T_2993 = ~ x3208_sm_io_output_ctr_inc;
  assign _T_3002 = x3208_sm_io_output_ctr_inc & _T_2996;
  assign _T_3009 = retime_released ? _T_3007 : 1'h0;
  assign _T_3018 = retime_released ? _T_3016 : 1'h0;
  assign _T_3025 = retime_released ? io_memStreams_loads_0_cmd_ready : 1'h0;
  assign _T_3026 = x3175_data_options_0[63:0];
  assign _T_3027 = x3175_data_options_0[95:64];
  assign _T_3028 = x3175_data_options_0[96];
  assign _T_3029 = ~ _T_3028;
  assign _T_3034 = retime_released ? x3177_now_valid : 1'h0;
  assign _T_3035 = x3236_en & retime_released;
  assign _T_3037 = x3236_sm_io_output_done;
  assign _T_3050 = retime_released ? _T_3048 : 1'h0;
  assign _T_3058 = retime_released ? _T_3056 : 1'h0;
  assign _T_3059 = ~ x3220_done;
  assign _T_3065 = retime_released ? _T_3063 : 1'h0;
  assign _T_3066 = _T_3058 & _T_3065;
  assign _T_3067 = ~ x3176_io_empty;
  assign _T_3073 = retime_released ? _T_3071 : 1'h0;
  assign _T_3075 = _T_3073 | _T_2886;
  assign _T_3076 = x3220_base_en & _T_3075;
  assign _T_3082 = retime_released ? _T_3080 : 1'h0;
  assign _T_3088 = retime_released ? _T_3086 : 1'h0;
  assign _T_3089 = ~ x3235_done;
  assign _T_3095 = retime_released ? _T_3093 : 1'h0;
  assign _T_3096 = _T_3088 & _T_3095;
  assign _T_3097 = x3235_base_en & x3177_valid;
  assign _T_3104 = x3220_en & retime_released;
  assign _T_3106 = x3220_sm_io_output_done;
  assign _T_3109 = x3220_sm_io_output_ctr_inc & _T_3059;
  assign _T_3110 = ~ x3220_ctr_trivial;
  assign _T_3111 = _T_3109 & _T_3110;
  assign _T_3112 = ~ x3220_sm_io_output_ctr_inc;
  assign _T_3121 = x3220_sm_io_output_ctr_inc & _T_3115;
  assign _T_3127 = retime_released ? _T_3125 : 1'h0;
  assign _T_3135 = retime_released ? _T_3133 : 1'h0;
  assign _T_3139 = $signed(x3221_number);
  assign _T_3408 = x3235_sm_io_output_done;
  assign _T_3410 = x3235_en & _T_3089;
  assign _T_3411 = ~ x3235_ctr_trivial;
  assign _T_3412 = _T_3410 & _T_3411;
  assign _T_3421 = retime_released ? _T_3419 : 1'h0;
  assign _T_3427 = retime_released ? _T_3425 : 1'h0;
  assign _T_3529 = $signed(_T_3504_number);
  assign _T_3530 = $signed(_T_3506_number);
  assign _T_3531 = $signed(_T_3529) < $signed(_T_3530);
  assign _T_3567 = retime_released ? _T_3565 : 1'h0;
  assign _T_3594 = _T_3569_number == 32'h0;
  assign _T_3595 = _T_3567 | _T_3594;
  assign _T_3596 = x3364_en & retime_released;
  assign _T_3598 = x3364_sm_io_output_done;
  assign _T_3611 = retime_released ? _T_3609 : 1'h0;
  assign _T_3619 = retime_released ? _T_3617 : 1'h0;
  assign _T_3620 = ~ x3335_done;
  assign _T_3626 = retime_released ? _T_3624 : 1'h0;
  assign _T_3627 = _T_3619 & _T_3626;
  assign _T_3628 = x3335_base_en & x3302_ready;
  assign _T_3629 = ~ x3303_io_full;
  assign _T_3635 = retime_released ? _T_3633 : 1'h0;
  assign _T_3636 = ~ b1204_chain_read_2;
  assign _T_3637 = _T_3635 | _T_3636;
  assign _T_3638 = _T_3628 & _T_3637;
  assign _T_3644 = retime_released ? _T_3642 : 1'h0;
  assign _T_3650 = retime_released ? _T_3648 : 1'h0;
  assign _T_3651 = ~ x3363_done;
  assign _T_3657 = retime_released ? _T_3655 : 1'h0;
  assign _T_3658 = _T_3650 & _T_3657;
  assign _T_3664 = retime_released ? _T_3662 : 1'h0;
  assign _T_3665 = x3427_en & retime_released;
  assign _T_3667 = x3427_sm_io_output_done;
  assign _T_3680 = retime_released ? _T_3678 : 1'h0;
  assign _T_3688 = retime_released ? _T_3686 : 1'h0;
  assign _T_3689 = ~ x3398_done;
  assign _T_3695 = retime_released ? _T_3693 : 1'h0;
  assign _T_3696 = _T_3688 & _T_3695;
  assign _T_3697 = x3398_base_en & x3365_ready;
  assign _T_3698 = ~ x3366_io_full;
  assign _T_3704 = retime_released ? _T_3702 : 1'h0;
  assign _T_3705 = ~ b1205_chain_read_2;
  assign _T_3706 = _T_3704 | _T_3705;
  assign _T_3707 = _T_3697 & _T_3706;
  assign _T_3713 = retime_released ? _T_3711 : 1'h0;
  assign _T_3719 = retime_released ? _T_3717 : 1'h0;
  assign _T_3720 = ~ x3426_done;
  assign _T_3726 = retime_released ? _T_3724 : 1'h0;
  assign _T_3727 = _T_3719 & _T_3726;
  assign _T_3733 = retime_released ? _T_3731 : 1'h0;
  assign _T_3734 = x3398_en & retime_released;
  assign _T_3736 = x3365_ready & _T_3698;
  assign _T_3737 = x3398_sm_io_output_done & _T_3736;
  assign _T_3740 = x3398_sm_io_output_ctr_inc & _T_3689;
  assign _T_3741 = ~ x3398_ctr_trivial;
  assign _T_3742 = _T_3740 & _T_3741;
  assign _T_3743 = ~ x3398_sm_io_output_ctr_inc;
  assign _T_3752 = x3398_sm_io_output_ctr_inc & _T_3746;
  assign _T_3759 = retime_released ? _T_3757 : 1'h0;
  assign _T_3768 = retime_released ? _T_3766 : 1'h0;
  assign _T_3775 = retime_released ? io_memStreams_loads_3_cmd_ready : 1'h0;
  assign _T_3776 = x3365_data_options_0[63:0];
  assign _T_3777 = x3365_data_options_0[95:64];
  assign _T_3778 = x3365_data_options_0[96];
  assign _T_3779 = ~ _T_3778;
  assign _T_3784 = retime_released ? x3367_now_valid : 1'h0;
  assign _T_3785 = x3426_en & retime_released;
  assign _T_3787 = x3426_sm_io_output_done;
  assign _T_3800 = retime_released ? _T_3798 : 1'h0;
  assign _T_3808 = retime_released ? _T_3806 : 1'h0;
  assign _T_3809 = ~ x3410_done;
  assign _T_3815 = retime_released ? _T_3813 : 1'h0;
  assign _T_3816 = _T_3808 & _T_3815;
  assign _T_3817 = ~ x3366_io_empty;
  assign _T_3823 = retime_released ? _T_3821 : 1'h0;
  assign _T_3825 = _T_3823 | _T_3705;
  assign _T_3826 = x3410_base_en & _T_3825;
  assign _T_3832 = retime_released ? _T_3830 : 1'h0;
  assign _T_3838 = retime_released ? _T_3836 : 1'h0;
  assign _T_3839 = ~ x3425_done;
  assign _T_3845 = retime_released ? _T_3843 : 1'h0;
  assign _T_3846 = _T_3838 & _T_3845;
  assign _T_3847 = x3425_base_en & x3367_valid;
  assign _GEN_0 = {{2'd0}, x3178_number};
  assign _T_3871 = _GEN_0 << 2;
  assign x3181 = x3179_number[5:0];
  assign _GEN_1 = {{2'd0}, x3183_number};
  assign _T_3874 = _GEN_1 << 2;
  assign _T_3891 = x3179_number[31];
  assign _T_3893 = {_T_3891,x3179_number};
  assign _T_3904 = x3182_number[31];
  assign _T_3906 = {_T_3904,x3182_number};
  assign _T_3907 = _T_3878_number - _T_3880_number;
  assign _T_3908 = $unsigned(_T_3907);
  assign _T_3909 = _T_3908[32:0];
  assign _T_3929 = _T_3876_number[31:0];
  assign _T_3959 = x3184_number[31];
  assign _T_3961 = {_T_3959,x3184_number};
  assign _T_3962 = _T_3933_number + _T_3935_number;
  assign _T_3963 = _T_3962[32:0];
  assign _T_3983 = _T_3931_number[31:0];
  assign x3188 = x3186_number[5:0];
  assign _T_4014 = _T_3989_number == 32'h0;
  assign _T_4048 = x3189_number[31];
  assign _T_4050 = {_T_4048,x3189_number};
  assign _T_4051 = 33'h40 - _T_4024_number;
  assign _T_4052 = $unsigned(_T_4051);
  assign _T_4053 = _T_4052[32:0];
  assign _T_4073 = _T_4020_number[31:0];
  assign _T_4078 = x3190 ? 32'h0 : x3191_number;
  assign _T_4085 = _T_3904 ? 2'h3 : 2'h0;
  assign _T_4086 = x3182_number[31:2];
  assign _T_4087 = {_T_4085,_T_4086};
  assign _T_4090 = x3192_number[31];
  assign _T_4094 = _T_4090 ? 2'h3 : 2'h0;
  assign _T_4095 = x3192_number[31:2];
  assign _T_4096 = {_T_4094,_T_4095};
  assign _T_4113 = x3193_number[31];
  assign _T_4115 = {_T_4113,x3193_number};
  assign _T_4126 = x3183_number[31];
  assign _T_4128 = {_T_4126,x3183_number};
  assign _T_4129 = _T_4100_number + _T_4102_number;
  assign _T_4130 = _T_4129[32:0];
  assign _T_4150 = _T_4098_number[31:0];
  assign _T_4183 = _T_4154_number + _T_4156_number;
  assign _T_4184 = _T_4183[32:0];
  assign _T_4204 = _T_4152_number[31:0];
  assign _T_4221 = x3196_number[31];
  assign _T_4223 = {_T_4221,x3196_number};
  assign _T_4234 = x3194_number[31];
  assign _T_4236 = {_T_4234,x3194_number};
  assign _T_4237 = _T_4208_number + _T_4210_number;
  assign _T_4238 = _T_4237[32:0];
  assign _T_4258 = _T_4206_number[31:0];
  assign _T_4291 = _T_4262_number + _T_4264_number;
  assign _T_4292 = _T_4291[32:0];
  assign _T_4312 = _T_4260_number[31:0];
  assign _T_4329 = x3198_number[31];
  assign _T_4331 = {_T_4329,x3198_number};
  assign _T_4344 = {_T_4090,x3192_number};
  assign _T_4345 = _T_4316_number + _T_4318_number;
  assign _T_4346 = _T_4345[32:0];
  assign _T_4366 = _T_4314_number[31:0];
  assign _T_4377 = x3185_number[31];
  assign _T_4381 = _T_4377 ? 32'hffffffff : 32'h0;
  assign _T_4383 = {_T_4381,x3185_number};
  assign _T_4415 = x3200_number[63];
  assign _T_4417 = {_T_4415,x3200_number};
  assign _T_4428 = _T_4385_number[63];
  assign _T_4430 = {_T_4428,_T_4385_number};
  assign _T_4431 = _T_4402_number + _T_4404_number;
  assign _T_4432 = _T_4431[64:0];
  assign _T_4452 = _T_4400_number[63:0];
  assign _T_4465 = {1'h1,x3204_item1};
  assign _T_4466 = {_T_4465,x3204_item0};
  assign _T_4472 = retime_released ? x3208_datapath_en : 1'h0;
  assign _T_4473 = _T_4472 & b1204_chain_read_1;
  assign _T_4480 = b1204_chain_read_1 & _T_4472;
  assign _T_4481 = {x3206_item2,x3206_item1};
  assign _T_4482 = {_T_4481,x3206_item0};
  assign _T_4503 = x3271_en & retime_released;
  assign _T_4505 = x3238_ready & _T_2948;
  assign _T_4506 = x3271_sm_io_output_done & _T_4505;
  assign _T_4509 = x3271_sm_io_output_ctr_inc & _T_2939;
  assign _T_4510 = ~ x3271_ctr_trivial;
  assign _T_4511 = _T_4509 & _T_4510;
  assign _T_4512 = ~ x3271_sm_io_output_ctr_inc;
  assign _T_4521 = x3271_sm_io_output_ctr_inc & _T_4515;
  assign _T_4528 = retime_released ? _T_4526 : 1'h0;
  assign _T_4537 = retime_released ? _T_4535 : 1'h0;
  assign _T_4544 = retime_released ? io_memStreams_loads_1_cmd_ready : 1'h0;
  assign _T_4545 = x3238_data_options_0[63:0];
  assign _T_4546 = x3238_data_options_0[95:64];
  assign _T_4547 = x3238_data_options_0[96];
  assign _T_4548 = ~ _T_4547;
  assign _T_4553 = retime_released ? x3240_now_valid : 1'h0;
  assign _T_4554 = x3299_en & retime_released;
  assign _T_4556 = x3299_sm_io_output_done;
  assign _T_4569 = retime_released ? _T_4567 : 1'h0;
  assign _T_4577 = retime_released ? _T_4575 : 1'h0;
  assign _T_4578 = ~ x3283_done;
  assign _T_4584 = retime_released ? _T_4582 : 1'h0;
  assign _T_4585 = _T_4577 & _T_4584;
  assign _T_4586 = ~ x3239_io_empty;
  assign _T_4592 = retime_released ? _T_4590 : 1'h0;
  assign _T_4594 = _T_4592 | _T_2955;
  assign _T_4595 = x3283_base_en & _T_4594;
  assign _T_4601 = retime_released ? _T_4599 : 1'h0;
  assign _T_4607 = retime_released ? _T_4605 : 1'h0;
  assign _T_4608 = ~ x3298_done;
  assign _T_4614 = retime_released ? _T_4612 : 1'h0;
  assign _T_4615 = _T_4607 & _T_4614;
  assign _T_4616 = x3298_base_en & x3240_valid;
  assign _T_4623 = x3283_en & retime_released;
  assign _T_4625 = x3283_sm_io_output_done;
  assign _T_4628 = x3283_sm_io_output_ctr_inc & _T_4578;
  assign _T_4629 = ~ x3283_ctr_trivial;
  assign _T_4630 = _T_4628 & _T_4629;
  assign _T_4631 = ~ x3283_sm_io_output_ctr_inc;
  assign _T_4640 = x3283_sm_io_output_ctr_inc & _T_4634;
  assign _T_4646 = retime_released ? _T_4644 : 1'h0;
  assign _T_4654 = retime_released ? _T_4652 : 1'h0;
  assign _T_4658 = $signed(x3284_number);
  assign _T_4927 = x3298_sm_io_output_done;
  assign _T_4929 = x3298_en & _T_4608;
  assign _T_4930 = ~ x3298_ctr_trivial;
  assign _T_4931 = _T_4929 & _T_4930;
  assign _T_4940 = retime_released ? _T_4938 : 1'h0;
  assign _T_4946 = retime_released ? _T_4944 : 1'h0;
  assign _T_5048 = $signed(_T_5023_number);
  assign _T_5049 = $signed(_T_5025_number);
  assign _T_5050 = $signed(_T_5048) < $signed(_T_5049);
  assign _T_5086 = retime_released ? _T_5084 : 1'h0;
  assign _T_5113 = _T_5088_number == 32'h0;
  assign _T_5114 = _T_5086 | _T_5113;
  assign _T_5115 = $signed(x3431_number);
  assign _T_5382 = x3466_en & retime_released;
  assign _T_5385 = retime_released ? x3466_sm_io_output_done : 1'h0;
  assign _T_5386 = ~ _T_5385;
  assign _T_5395 = _T_5385 & _T_5389;
  assign _T_5397 = x3466_sm_io_output_ctr_inc & _T_2764;
  assign _T_5398 = ~ x3466_ctr_trivial;
  assign _T_5399 = _T_5397 & _T_5398;
  assign _T_5400 = x3466_sm_io_output_ctr_inc;
  assign _T_5403 = retime_released ? x3466_rst_en : 1'h0;
  assign _T_5409 = retime_released ? _T_5407 : 1'h0;
  assign _T_5416 = x3466_datapath_en & _T_2764;
  assign _T_5516 = $signed(_T_5491_number);
  assign _T_5517 = $signed(_T_5493_number);
  assign _T_5518 = $signed(_T_5516) < $signed(_T_5517);
  assign _T_5646 = $signed(_T_5621_number);
  assign _T_5647 = $signed(_T_5623_number);
  assign _T_5648 = $signed(_T_5646) < $signed(_T_5647);
  assign _T_5776 = $signed(_T_5751_number);
  assign _T_5777 = $signed(_T_5753_number);
  assign _T_5778 = $signed(_T_5776) < $signed(_T_5777);
  assign _T_5906 = $signed(_T_5881_number);
  assign _T_5907 = $signed(_T_5883_number);
  assign _T_5908 = $signed(_T_5906) < $signed(_T_5907);
  assign _T_5944 = retime_released ? _T_5942 : 1'h0;
  assign _T_5971 = _T_5946_number == 32'h0;
  assign _T_5972 = _T_5944 | _T_5971;
  assign _T_5973 = $signed(x3467_number);
  assign _T_6240 = x3502_en & retime_released;
  assign _T_6243 = retime_released ? x3502_sm_io_output_done : 1'h0;
  assign _T_6244 = ~ _T_6243;
  assign _T_6253 = _T_6243 & _T_6247;
  assign _T_6255 = x3502_sm_io_output_ctr_inc & _T_2784;
  assign _T_6256 = ~ x3502_ctr_trivial;
  assign _T_6257 = _T_6255 & _T_6256;
  assign _T_6258 = x3502_sm_io_output_ctr_inc;
  assign _T_6261 = retime_released ? x3502_rst_en : 1'h0;
  assign _T_6267 = retime_released ? _T_6265 : 1'h0;
  assign _T_6274 = x3502_datapath_en & _T_2784;
  assign _T_6374 = $signed(_T_6349_number);
  assign _T_6375 = $signed(_T_6351_number);
  assign _T_6376 = $signed(_T_6374) < $signed(_T_6375);
  assign _T_6504 = $signed(_T_6479_number);
  assign _T_6505 = $signed(_T_6481_number);
  assign _T_6506 = $signed(_T_6504) < $signed(_T_6505);
  assign _T_6634 = $signed(_T_6609_number);
  assign _T_6635 = $signed(_T_6611_number);
  assign _T_6636 = $signed(_T_6634) < $signed(_T_6635);
  assign _T_6764 = $signed(_T_6739_number);
  assign _T_6765 = $signed(_T_6741_number);
  assign _T_6766 = $signed(_T_6764) < $signed(_T_6765);
  assign _T_6802 = retime_released ? _T_6800 : 1'h0;
  assign _T_6829 = _T_6804_number == 32'h0;
  assign _T_6830 = _T_6802 | _T_6829;
  assign _T_6845 = x3505_number[7:0];
  assign _T_6846 = x3505_number[31];
  assign _T_6847 = x3505_number[31:8];
  assign _T_6848 = {_T_6846,_T_6847};
  assign _T_6849 = {_T_6844,_T_6842};
  assign _T_6858 = x3504_number[7:0];
  assign _T_6859 = x3504_number[31];
  assign _T_6860 = x3504_number[31:8];
  assign _T_6861 = {_T_6859,_T_6860};
  assign _T_6862 = {_T_6857,_T_6855};
  assign _T_6863 = _T_6834_number + _T_6836_number;
  assign _T_6864 = _T_6863[32:0];
  assign _T_6881 = _T_6832_number[7:0];
  assign _T_6883 = _T_6832_number[31:8];
  assign _T_6884 = {_T_6880,_T_6878};
  assign _T_6885 = b1205_chain_read_4 ? x3506_number : x3505_number;
  assign _T_6934 = _T_6909_number == 32'h0;
  assign _T_6949 = x3507_number[7:0];
  assign _T_6950 = x3507_number[31];
  assign _T_6951 = x3507_number[31:8];
  assign _T_6952 = {_T_6950,_T_6951};
  assign _T_6953 = {_T_6948,_T_6946};
  assign _T_6967 = _T_6938_number + 33'h0;
  assign _T_6968 = _T_6967[32:0];
  assign _T_6985 = _T_6936_number[7:0];
  assign _T_6987 = _T_6936_number[31:8];
  assign _T_6988 = {_T_6984,_T_6982};
  assign _T_6989 = x3510 ? x3507_number : x3511_number;
  assign _T_6997 = retime_released ? _T_6995 : 1'h0;
  assign _T_7005 = retime_released ? x3152_wren : 1'h0;
  assign _T_7008 = retime_released ? x3152_resetter : 1'h0;
  assign _T_7009 = reset | _T_7008;
  assign _T_7010 = x3516_number[31];
  assign _T_7014 = _T_7010 ? 32'hffffffff : 32'h0;
  assign _T_7015 = {_T_7014,x3516_number};
  assign _GEN_2 = {{2'd0}, x3241_number};
  assign _T_7036 = _GEN_2 << 2;
  assign x3244 = x3242_number[5:0];
  assign _GEN_3 = {{2'd0}, x3246_number};
  assign _T_7039 = _GEN_3 << 2;
  assign _T_7056 = x3242_number[31];
  assign _T_7058 = {_T_7056,x3242_number};
  assign _T_7069 = x3245_number[31];
  assign _T_7071 = {_T_7069,x3245_number};
  assign _T_7072 = _T_7043_number - _T_7045_number;
  assign _T_7073 = $unsigned(_T_7072);
  assign _T_7074 = _T_7073[32:0];
  assign _T_7094 = _T_7041_number[31:0];
  assign _T_7124 = x3247_number[31];
  assign _T_7126 = {_T_7124,x3247_number};
  assign _T_7127 = _T_7098_number + _T_7100_number;
  assign _T_7128 = _T_7127[32:0];
  assign _T_7148 = _T_7096_number[31:0];
  assign x3251 = x3249_number[5:0];
  assign _T_7179 = _T_7154_number == 32'h0;
  assign _T_7213 = x3252_number[31];
  assign _T_7215 = {_T_7213,x3252_number};
  assign _T_7216 = 33'h40 - _T_7189_number;
  assign _T_7217 = $unsigned(_T_7216);
  assign _T_7218 = _T_7217[32:0];
  assign _T_7238 = _T_7185_number[31:0];
  assign _T_7243 = x3253 ? 32'h0 : x3254_number;
  assign _T_7250 = _T_7069 ? 2'h3 : 2'h0;
  assign _T_7251 = x3245_number[31:2];
  assign _T_7252 = {_T_7250,_T_7251};
  assign _T_7255 = x3255_number[31];
  assign _T_7259 = _T_7255 ? 2'h3 : 2'h0;
  assign _T_7260 = x3255_number[31:2];
  assign _T_7261 = {_T_7259,_T_7260};
  assign _T_7278 = x3256_number[31];
  assign _T_7280 = {_T_7278,x3256_number};
  assign _T_7291 = x3246_number[31];
  assign _T_7293 = {_T_7291,x3246_number};
  assign _T_7294 = _T_7265_number + _T_7267_number;
  assign _T_7295 = _T_7294[32:0];
  assign _T_7315 = _T_7263_number[31:0];
  assign _T_7348 = _T_7319_number + _T_7321_number;
  assign _T_7349 = _T_7348[32:0];
  assign _T_7369 = _T_7317_number[31:0];
  assign _T_7386 = x3259_number[31];
  assign _T_7388 = {_T_7386,x3259_number};
  assign _T_7399 = x3257_number[31];
  assign _T_7401 = {_T_7399,x3257_number};
  assign _T_7402 = _T_7373_number + _T_7375_number;
  assign _T_7403 = _T_7402[32:0];
  assign _T_7423 = _T_7371_number[31:0];
  assign _T_7456 = _T_7427_number + _T_7429_number;
  assign _T_7457 = _T_7456[32:0];
  assign _T_7477 = _T_7425_number[31:0];
  assign _T_7494 = x3261_number[31];
  assign _T_7496 = {_T_7494,x3261_number};
  assign _T_7509 = {_T_7255,x3255_number};
  assign _T_7510 = _T_7481_number + _T_7483_number;
  assign _T_7511 = _T_7510[32:0];
  assign _T_7531 = _T_7479_number[31:0];
  assign _T_7542 = x3248_number[31];
  assign _T_7546 = _T_7542 ? 32'hffffffff : 32'h0;
  assign _T_7548 = {_T_7546,x3248_number};
  assign _T_7580 = x3263_number[63];
  assign _T_7582 = {_T_7580,x3263_number};
  assign _T_7593 = _T_7550_number[63];
  assign _T_7595 = {_T_7593,_T_7550_number};
  assign _T_7596 = _T_7567_number + _T_7569_number;
  assign _T_7597 = _T_7596[64:0];
  assign _T_7617 = _T_7565_number[63:0];
  assign _T_7630 = {1'h1,x3267_item1};
  assign _T_7631 = {_T_7630,x3267_item0};
  assign _T_7637 = retime_released ? x3271_datapath_en : 1'h0;
  assign _T_7638 = _T_7637 & b1205_chain_read_1;
  assign _T_7645 = b1205_chain_read_1 & _T_7637;
  assign _T_7646 = {x3269_item2,x3269_item1};
  assign _T_7647 = {_T_7646,x3269_item0};
  assign _GEN_4 = {{2'd0}, x3368_number};
  assign _T_7685 = _GEN_4 << 2;
  assign x3371 = x3369_number[5:0];
  assign _GEN_5 = {{2'd0}, x3373_number};
  assign _T_7688 = _GEN_5 << 2;
  assign _T_7705 = x3369_number[31];
  assign _T_7707 = {_T_7705,x3369_number};
  assign _T_7718 = x3372_number[31];
  assign _T_7720 = {_T_7718,x3372_number};
  assign _T_7721 = _T_7692_number - _T_7694_number;
  assign _T_7722 = $unsigned(_T_7721);
  assign _T_7723 = _T_7722[32:0];
  assign _T_7743 = _T_7690_number[31:0];
  assign _T_7773 = x3374_number[31];
  assign _T_7775 = {_T_7773,x3374_number};
  assign _T_7776 = _T_7747_number + _T_7749_number;
  assign _T_7777 = _T_7776[32:0];
  assign _T_7797 = _T_7745_number[31:0];
  assign x3378 = x3376_number[5:0];
  assign _T_7828 = _T_7803_number == 32'h0;
  assign _T_7862 = x3379_number[31];
  assign _T_7864 = {_T_7862,x3379_number};
  assign _T_7865 = 33'h40 - _T_7838_number;
  assign _T_7866 = $unsigned(_T_7865);
  assign _T_7867 = _T_7866[32:0];
  assign _T_7887 = _T_7834_number[31:0];
  assign _T_7892 = x3380 ? 32'h0 : x3381_number;
  assign _T_7899 = _T_7718 ? 2'h3 : 2'h0;
  assign _T_7900 = x3372_number[31:2];
  assign _T_7901 = {_T_7899,_T_7900};
  assign _T_7904 = x3382_number[31];
  assign _T_7908 = _T_7904 ? 2'h3 : 2'h0;
  assign _T_7909 = x3382_number[31:2];
  assign _T_7910 = {_T_7908,_T_7909};
  assign _T_7927 = x3383_number[31];
  assign _T_7929 = {_T_7927,x3383_number};
  assign _T_7940 = x3373_number[31];
  assign _T_7942 = {_T_7940,x3373_number};
  assign _T_7943 = _T_7914_number + _T_7916_number;
  assign _T_7944 = _T_7943[32:0];
  assign _T_7964 = _T_7912_number[31:0];
  assign _T_7997 = _T_7968_number + _T_7970_number;
  assign _T_7998 = _T_7997[32:0];
  assign _T_8018 = _T_7966_number[31:0];
  assign _T_8035 = x3386_number[31];
  assign _T_8037 = {_T_8035,x3386_number};
  assign _T_8048 = x3384_number[31];
  assign _T_8050 = {_T_8048,x3384_number};
  assign _T_8051 = _T_8022_number + _T_8024_number;
  assign _T_8052 = _T_8051[32:0];
  assign _T_8072 = _T_8020_number[31:0];
  assign _T_8105 = _T_8076_number + _T_8078_number;
  assign _T_8106 = _T_8105[32:0];
  assign _T_8126 = _T_8074_number[31:0];
  assign _T_8143 = x3388_number[31];
  assign _T_8145 = {_T_8143,x3388_number};
  assign _T_8158 = {_T_7904,x3382_number};
  assign _T_8159 = _T_8130_number + _T_8132_number;
  assign _T_8160 = _T_8159[32:0];
  assign _T_8180 = _T_8128_number[31:0];
  assign _T_8191 = x3375_number[31];
  assign _T_8195 = _T_8191 ? 32'hffffffff : 32'h0;
  assign _T_8197 = {_T_8195,x3375_number};
  assign _T_8229 = x3390_number[63];
  assign _T_8231 = {_T_8229,x3390_number};
  assign _T_8242 = _T_8199_number[63];
  assign _T_8244 = {_T_8242,_T_8199_number};
  assign _T_8245 = _T_8216_number + _T_8218_number;
  assign _T_8246 = _T_8245[64:0];
  assign _T_8266 = _T_8214_number[63:0];
  assign _T_8279 = {1'h1,x3394_item1};
  assign _T_8280 = {_T_8279,x3394_item0};
  assign _T_8286 = retime_released ? x3398_datapath_en : 1'h0;
  assign _T_8287 = _T_8286 & b1205_chain_read_2;
  assign _T_8294 = b1205_chain_read_2 & _T_8286;
  assign _T_8295 = {x3396_item2,x3396_item1};
  assign _T_8296 = {_T_8295,x3396_item0};
  assign _T_8317 = x3167_en & retime_released;
  assign _T_8320 = retime_released ? x3167_sm_io_output_done : 1'h0;
  assign _T_8321 = ~ _T_8320;
  assign _T_8330 = _T_8320 & _T_8324;
  assign _T_8333 = x3167_sm_io_output_ctr_inc & _T_2552;
  assign _T_8334 = ~ x3167_ctr_trivial;
  assign _T_8335 = _T_8333 & _T_8334;
  assign _T_8336 = ~ x3167_sm_io_output_ctr_inc;
  assign _T_8345 = x3167_sm_io_output_ctr_inc & _T_8339;
  assign _T_8351 = retime_released ? _T_8349 : 1'h0;
  assign _T_8359 = retime_released ? _T_8357 : 1'h0;
  assign _T_8363 = x3173_en & retime_released;
  assign _T_8366 = retime_released ? x3173_sm_io_output_done : 1'h0;
  assign _T_8367 = ~ _T_8366;
  assign _T_8376 = _T_8366 & _T_8370;
  assign _T_8379 = x3173_sm_io_output_ctr_inc & _T_2572;
  assign _T_8380 = ~ x3173_ctr_trivial;
  assign _T_8381 = _T_8379 & _T_8380;
  assign _T_8382 = ~ x3173_sm_io_output_ctr_inc;
  assign _T_8391 = x3173_sm_io_output_ctr_inc & _T_8385;
  assign _T_8397 = retime_released ? _T_8395 : 1'h0;
  assign _T_8405 = retime_released ? _T_8403 : 1'h0;
  assign _T_8425 = x3168_number[31];
  assign _T_8427 = {_T_8425,x3168_number};
  assign _T_8438 = b1203_number[31];
  assign _T_8440 = {_T_8438,b1203_number};
  assign _T_8441 = _T_8412_number - _T_8414_number;
  assign _T_8442 = $unsigned(_T_8441);
  assign _T_8443 = _T_8442[32:0];
  assign _T_8463 = _T_8410_number[31:0];
  assign _T_8495 = $signed(_T_8471_number);
  assign _T_8496 = $signed(32'sh40) < $signed(_T_8495);
  assign _T_8501_number = _T_8496 ? 32'h40 : x3169_number;
  assign _T_8559 = retime_released ? x3173_datapath_en : 1'h0;
  assign _T_8560 = b1205 & _T_8559;
  assign _T_8565 = ~ _T_8560;
  assign _T_8566 = _T_8564 & _T_8565;
  assign _T_8573 = retime_released ? _T_8571 : 1'h0;
  assign _T_8579 = retime_released ? _T_8577 : 1'h0;
  assign _T_8585 = retime_released ? _T_8583 : 1'h0;
  assign _T_8591 = retime_released ? _T_8589 : 1'h0;
  assign _T_8597 = retime_released ? _T_8595 : 1'h0;
  assign _T_8603 = retime_released ? _T_8601 : 1'h0;
  assign _T_8609 = retime_released ? _T_8607 : 1'h0;
  assign _T_8615 = retime_released ? _T_8613 : 1'h0;
  assign _T_8621 = retime_released ? _T_8619 : 1'h0;
  assign _T_8627 = retime_released ? _T_8625 : 1'h0;
  assign _T_8630 = retime_released ? x3174_done : 1'h0;
  assign _T_8633 = retime_released ? x3301_done : 1'h0;
  assign _T_8636 = retime_released ? x3428_done : 1'h0;
  assign _T_8639 = retime_released ? x3503_done : 1'h0;
  assign _T_8642 = retime_released ? x3514_done : 1'h0;
  assign _T_8663 = retime_released ? _T_8661 : 1'h0;
  assign _T_8669 = retime_released ? _T_8667 : 1'h0;
  assign _T_8675 = retime_released ? _T_8673 : 1'h0;
  assign _T_8681 = retime_released ? _T_8679 : 1'h0;
  assign _T_8687 = retime_released ? _T_8685 : 1'h0;
  assign _T_8693 = retime_released ? _T_8691 : 1'h0;
  assign _T_8699 = retime_released ? _T_8697 : 1'h0;
  assign _T_8705 = retime_released ? _T_8703 : 1'h0;
  assign _T_8711 = retime_released ? _T_8709 : 1'h0;
  assign _T_8717 = retime_released ? _T_8715 : 1'h0;
  assign _T_8723 = retime_released ? _T_8721 : 1'h0;
  assign _T_8729 = retime_released ? _T_8727 : 1'h0;
  assign _T_8735 = retime_released ? _T_8733 : 1'h0;
  assign _T_8741 = retime_released ? _T_8739 : 1'h0;
  assign _T_8747 = retime_released ? _T_8745 : 1'h0;
  assign _T_8753 = retime_released ? _T_8751 : 1'h0;
  assign _T_8759 = retime_released ? _T_8757 : 1'h0;
  assign _T_8765 = retime_released ? _T_8763 : 1'h0;
  assign _T_8771 = retime_released ? _T_8769 : 1'h0;
  assign _T_8777 = retime_released ? _T_8775 : 1'h0;
  assign _T_8783 = retime_released ? _T_8781 : 1'h0;
  assign _T_8789 = retime_released ? _T_8787 : 1'h0;
  assign _T_8790 = $unsigned(x3468_0);
  assign _T_8791 = $unsigned(x3468_1);
  assign _T_8792 = $unsigned(x3468_2);
  assign _T_8793 = $unsigned(x3468_3);
  assign _T_8794 = b1524 & b1205_chain_read_3;
  assign _T_8795 = b1525 & b1205_chain_read_3;
  assign _T_8796 = b1526 & b1205_chain_read_3;
  assign _T_8797 = b1527 & b1205_chain_read_3;
  assign _T_8800 = retime_released ? x3502_en : 1'h0;
  assign _T_8801 = _T_8800 & x3470;
  assign _T_8805 = _T_8800 & x3471;
  assign _T_8809 = _T_8800 & x3472;
  assign _T_8813 = _T_8800 & x3473;
  assign _T_8900 = x3475_number[31];
  assign _T_8904 = _T_8900 ? 8'hff : 8'h0;
  assign _T_8905 = {_T_8904,x3475_number};
  assign _T_8906 = x3480_number[31];
  assign _T_8910 = _T_8906 ? 8'hff : 8'h0;
  assign _T_8911 = {_T_8910,x3480_number};
  assign _T_8912 = _T_8905 * _T_8911;
  assign _T_8913 = _T_8912[79:8];
  assign _T_8931 = _T_8899_number[7:0];
  assign _T_8932 = _T_8899_number[31:8];
  assign _T_8933 = {_T_8930,_T_8928};
  assign _T_8936 = x3476_number[31];
  assign _T_8940 = _T_8936 ? 8'hff : 8'h0;
  assign _T_8941 = {_T_8940,x3476_number};
  assign _T_8942 = x3481_number[31];
  assign _T_8946 = _T_8942 ? 8'hff : 8'h0;
  assign _T_8947 = {_T_8946,x3481_number};
  assign _T_8948 = _T_8941 * _T_8947;
  assign _T_8949 = _T_8948[79:8];
  assign _T_8967 = _T_8935_number[7:0];
  assign _T_8968 = _T_8935_number[31:8];
  assign _T_8969 = {_T_8966,_T_8964};
  assign _T_8972 = x3477_number[31];
  assign _T_8976 = _T_8972 ? 8'hff : 8'h0;
  assign _T_8977 = {_T_8976,x3477_number};
  assign _T_8978 = x3482_number[31];
  assign _T_8982 = _T_8978 ? 8'hff : 8'h0;
  assign _T_8983 = {_T_8982,x3482_number};
  assign _T_8984 = _T_8977 * _T_8983;
  assign _T_8985 = _T_8984[79:8];
  assign _T_9003 = _T_8971_number[7:0];
  assign _T_9004 = _T_8971_number[31:8];
  assign _T_9005 = {_T_9002,_T_9000};
  assign _T_9008 = x3478_number[31];
  assign _T_9012 = _T_9008 ? 8'hff : 8'h0;
  assign _T_9013 = {_T_9012,x3478_number};
  assign _T_9014 = x3483_number[31];
  assign _T_9018 = _T_9014 ? 8'hff : 8'h0;
  assign _T_9019 = {_T_9018,x3483_number};
  assign _T_9020 = _T_9013 * _T_9019;
  assign _T_9021 = _T_9020[79:8];
  assign _T_9039 = _T_9007_number[7:0];
  assign _T_9040 = _T_9007_number[31:8];
  assign _T_9041 = {_T_9038,_T_9036};
  assign _T_9056 = x3484_number[7:0];
  assign _T_9057 = x3484_number[31];
  assign _T_9058 = x3484_number[31:8];
  assign _T_9059 = {_T_9057,_T_9058};
  assign _T_9060 = {_T_9055,_T_9053};
  assign _T_9069 = x3485_number[7:0];
  assign _T_9070 = x3485_number[31];
  assign _T_9071 = x3485_number[31:8];
  assign _T_9072 = {_T_9070,_T_9071};
  assign _T_9073 = {_T_9068,_T_9066};
  assign _T_9074 = _T_9045_number + _T_9047_number;
  assign _T_9075 = _T_9074[32:0];
  assign _T_9092 = _T_9043_number[7:0];
  assign _T_9094 = _T_9043_number[31:8];
  assign _T_9095 = {_T_9091,_T_9089};
  assign _T_9096 = x3471 ? x3488_number : x3484_number;
  assign _T_9112 = x3486_number[7:0];
  assign _T_9113 = x3486_number[31];
  assign _T_9114 = x3486_number[31:8];
  assign _T_9115 = {_T_9113,_T_9114};
  assign _T_9116 = {_T_9111,_T_9109};
  assign _T_9125 = x3487_number[7:0];
  assign _T_9126 = x3487_number[31];
  assign _T_9127 = x3487_number[31:8];
  assign _T_9128 = {_T_9126,_T_9127};
  assign _T_9129 = {_T_9124,_T_9122};
  assign _T_9130 = _T_9101_number + _T_9103_number;
  assign _T_9131 = _T_9130[32:0];
  assign _T_9148 = _T_9099_number[7:0];
  assign _T_9150 = _T_9099_number[31:8];
  assign _T_9151 = {_T_9147,_T_9145};
  assign _T_9152 = x3473 ? x3491_number : x3486_number;
  assign _T_9153 = x3472 | x3473;
  assign _T_9168 = x3489_number[7:0];
  assign _T_9169 = x3489_number[31];
  assign _T_9170 = x3489_number[31:8];
  assign _T_9171 = {_T_9169,_T_9170};
  assign _T_9172 = {_T_9167,_T_9165};
  assign _T_9181 = x3492_number[7:0];
  assign _T_9182 = x3492_number[31];
  assign _T_9183 = x3492_number[31:8];
  assign _T_9184 = {_T_9182,_T_9183};
  assign _T_9185 = {_T_9180,_T_9178};
  assign _T_9186 = _T_9157_number + _T_9159_number;
  assign _T_9187 = _T_9186[32:0];
  assign _T_9204 = _T_9155_number[7:0];
  assign _T_9206 = _T_9155_number[31:8];
  assign _T_9207 = {_T_9203,_T_9201};
  assign _T_9208 = x3493 ? x3494_number : x3489_number;
  assign _T_9242 = _T_9217_number == 32'h0;
  assign _T_9257 = x3495_number[7:0];
  assign _T_9258 = x3495_number[31];
  assign _T_9259 = x3495_number[31:8];
  assign _T_9260 = {_T_9258,_T_9259};
  assign _T_9261 = {_T_9256,_T_9254};
  assign _T_9275 = _T_9246_number + 33'h0;
  assign _T_9276 = _T_9275[32:0];
  assign _T_9293 = _T_9244_number[7:0];
  assign _T_9295 = _T_9244_number[31:8];
  assign _T_9296 = {_T_9292,_T_9290};
  assign _T_9297 = x3498 ? x3495_number : x3499_number;
  assign _T_9300 = retime_released ? x3430_wren : 1'h0;
  assign _T_9303 = retime_released ? x3430_resetter : 1'h0;
  assign _T_9304 = reset | _T_9303;
  assign _T_9311 = retime_released ? _T_9309 : 1'h0;
  assign _T_9312 = b1205_chain_read_3 & _T_9311;
  assign _T_9318 = x3335_en & retime_released;
  assign _T_9320 = x3302_ready & _T_3629;
  assign _T_9321 = x3335_sm_io_output_done & _T_9320;
  assign _T_9324 = x3335_sm_io_output_ctr_inc & _T_3620;
  assign _T_9325 = ~ x3335_ctr_trivial;
  assign _T_9326 = _T_9324 & _T_9325;
  assign _T_9327 = ~ x3335_sm_io_output_ctr_inc;
  assign _T_9336 = x3335_sm_io_output_ctr_inc & _T_9330;
  assign _T_9343 = retime_released ? _T_9341 : 1'h0;
  assign _T_9352 = retime_released ? _T_9350 : 1'h0;
  assign _T_9359 = retime_released ? io_memStreams_loads_2_cmd_ready : 1'h0;
  assign _T_9360 = x3302_data_options_0[63:0];
  assign _T_9361 = x3302_data_options_0[95:64];
  assign _T_9362 = x3302_data_options_0[96];
  assign _T_9363 = ~ _T_9362;
  assign _T_9368 = retime_released ? x3304_now_valid : 1'h0;
  assign _T_9369 = x3363_en & retime_released;
  assign _T_9371 = x3363_sm_io_output_done;
  assign _T_9384 = retime_released ? _T_9382 : 1'h0;
  assign _T_9392 = retime_released ? _T_9390 : 1'h0;
  assign _T_9393 = ~ x3347_done;
  assign _T_9399 = retime_released ? _T_9397 : 1'h0;
  assign _T_9400 = _T_9392 & _T_9399;
  assign _T_9401 = ~ x3303_io_empty;
  assign _T_9407 = retime_released ? _T_9405 : 1'h0;
  assign _T_9409 = _T_9407 | _T_3636;
  assign _T_9410 = x3347_base_en & _T_9409;
  assign _T_9416 = retime_released ? _T_9414 : 1'h0;
  assign _T_9422 = retime_released ? _T_9420 : 1'h0;
  assign _T_9423 = ~ x3362_done;
  assign _T_9429 = retime_released ? _T_9427 : 1'h0;
  assign _T_9430 = _T_9422 & _T_9429;
  assign _T_9431 = x3362_base_en & x3304_valid;
  assign _T_9438 = x3347_en & retime_released;
  assign _T_9440 = x3347_sm_io_output_done;
  assign _T_9443 = x3347_sm_io_output_ctr_inc & _T_9393;
  assign _T_9444 = ~ x3347_ctr_trivial;
  assign _T_9445 = _T_9443 & _T_9444;
  assign _T_9446 = ~ x3347_sm_io_output_ctr_inc;
  assign _T_9455 = x3347_sm_io_output_ctr_inc & _T_9449;
  assign _T_9461 = retime_released ? _T_9459 : 1'h0;
  assign _T_9469 = retime_released ? _T_9467 : 1'h0;
  assign _T_9473 = $signed(x3348_number);
  assign _T_9742 = x3362_sm_io_output_done;
  assign _T_9744 = x3362_en & _T_9423;
  assign _T_9745 = ~ x3362_ctr_trivial;
  assign _T_9746 = _T_9744 & _T_9745;
  assign _T_9755 = retime_released ? _T_9753 : 1'h0;
  assign _T_9761 = retime_released ? _T_9759 : 1'h0;
  assign _T_9863 = $signed(_T_9838_number);
  assign _T_9864 = $signed(_T_9840_number);
  assign _T_9865 = $signed(_T_9863) < $signed(_T_9864);
  assign _T_9901 = retime_released ? _T_9899 : 1'h0;
  assign _T_9928 = _T_9903_number == 32'h0;
  assign _T_9929 = _T_9901 | _T_9928;
  assign _T_9930 = $unsigned(x3349_0);
  assign _T_9957 = $signed(_T_9932_number);
  assign _T_9958 = $signed(_T_9934_number);
  assign _T_9959 = $signed(_T_9957) <= $signed(_T_9958);
  assign _T_9986 = $signed(_T_9961_number);
  assign _T_9987 = $signed(_T_9963_number);
  assign _T_9988 = $signed(_T_9986) < $signed(_T_9987);
  assign _T_9989 = x3352 & x3354;
  assign _T_10006 = b1393_number[31];
  assign _T_10008 = {_T_10006,b1393_number};
  assign _T_10019 = x3351_number[31];
  assign _T_10021 = {_T_10019,x3351_number};
  assign _T_10022 = _T_9993_number - _T_9995_number;
  assign _T_10023 = $unsigned(_T_10022);
  assign _T_10024 = _T_10023[32:0];
  assign _T_10044 = _T_9991_number[31:0];
  assign _T_10045 = b1394 & b1204_chain_read_2;
  assign _T_10048 = x3357 & x3362_datapath_en;
  assign _T_10049 = x3355 & x3357;
  assign _T_10054 = x3360 & x3362_datapath_en;
  assign _T_10055 = $unsigned(x3432_0);
  assign _T_10056 = $unsigned(x3432_1);
  assign _T_10057 = $unsigned(x3432_2);
  assign _T_10058 = $unsigned(x3432_3);
  assign _T_10059 = b1483 & b1204_chain_read_3;
  assign _T_10060 = b1484 & b1204_chain_read_3;
  assign _T_10061 = b1485 & b1204_chain_read_3;
  assign _T_10062 = b1486 & b1204_chain_read_3;
  assign _T_10065 = retime_released ? x3466_en : 1'h0;
  assign _T_10066 = _T_10065 & x3434;
  assign _T_10070 = _T_10065 & x3435;
  assign _T_10074 = _T_10065 & x3436;
  assign _T_10078 = _T_10065 & x3437;
  assign _T_10165 = x3439_number[31];
  assign _T_10169 = _T_10165 ? 8'hff : 8'h0;
  assign _T_10170 = {_T_10169,x3439_number};
  assign _T_10171 = x3444_number[31];
  assign _T_10175 = _T_10171 ? 8'hff : 8'h0;
  assign _T_10176 = {_T_10175,x3444_number};
  assign _T_10177 = _T_10170 * _T_10176;
  assign _T_10178 = _T_10177[79:8];
  assign _T_10196 = _T_10164_number[7:0];
  assign _T_10197 = _T_10164_number[31:8];
  assign _T_10198 = {_T_10195,_T_10193};
  assign _T_10201 = x3440_number[31];
  assign _T_10205 = _T_10201 ? 8'hff : 8'h0;
  assign _T_10206 = {_T_10205,x3440_number};
  assign _T_10207 = x3445_number[31];
  assign _T_10211 = _T_10207 ? 8'hff : 8'h0;
  assign _T_10212 = {_T_10211,x3445_number};
  assign _T_10213 = _T_10206 * _T_10212;
  assign _T_10214 = _T_10213[79:8];
  assign _T_10232 = _T_10200_number[7:0];
  assign _T_10233 = _T_10200_number[31:8];
  assign _T_10234 = {_T_10231,_T_10229};
  assign _T_10237 = x3441_number[31];
  assign _T_10241 = _T_10237 ? 8'hff : 8'h0;
  assign _T_10242 = {_T_10241,x3441_number};
  assign _T_10243 = x3446_number[31];
  assign _T_10247 = _T_10243 ? 8'hff : 8'h0;
  assign _T_10248 = {_T_10247,x3446_number};
  assign _T_10249 = _T_10242 * _T_10248;
  assign _T_10250 = _T_10249[79:8];
  assign _T_10268 = _T_10236_number[7:0];
  assign _T_10269 = _T_10236_number[31:8];
  assign _T_10270 = {_T_10267,_T_10265};
  assign _T_10273 = x3442_number[31];
  assign _T_10277 = _T_10273 ? 8'hff : 8'h0;
  assign _T_10278 = {_T_10277,x3442_number};
  assign _T_10279 = x3447_number[31];
  assign _T_10283 = _T_10279 ? 8'hff : 8'h0;
  assign _T_10284 = {_T_10283,x3447_number};
  assign _T_10285 = _T_10278 * _T_10284;
  assign _T_10286 = _T_10285[79:8];
  assign _T_10304 = _T_10272_number[7:0];
  assign _T_10305 = _T_10272_number[31:8];
  assign _T_10306 = {_T_10303,_T_10301};
  assign _T_10321 = x3448_number[7:0];
  assign _T_10322 = x3448_number[31];
  assign _T_10323 = x3448_number[31:8];
  assign _T_10324 = {_T_10322,_T_10323};
  assign _T_10325 = {_T_10320,_T_10318};
  assign _T_10334 = x3449_number[7:0];
  assign _T_10335 = x3449_number[31];
  assign _T_10336 = x3449_number[31:8];
  assign _T_10337 = {_T_10335,_T_10336};
  assign _T_10338 = {_T_10333,_T_10331};
  assign _T_10339 = _T_10310_number + _T_10312_number;
  assign _T_10340 = _T_10339[32:0];
  assign _T_10357 = _T_10308_number[7:0];
  assign _T_10359 = _T_10308_number[31:8];
  assign _T_10360 = {_T_10356,_T_10354};
  assign _T_10361 = x3435 ? x3452_number : x3448_number;
  assign _T_10377 = x3450_number[7:0];
  assign _T_10378 = x3450_number[31];
  assign _T_10379 = x3450_number[31:8];
  assign _T_10380 = {_T_10378,_T_10379};
  assign _T_10381 = {_T_10376,_T_10374};
  assign _T_10390 = x3451_number[7:0];
  assign _T_10391 = x3451_number[31];
  assign _T_10392 = x3451_number[31:8];
  assign _T_10393 = {_T_10391,_T_10392};
  assign _T_10394 = {_T_10389,_T_10387};
  assign _T_10395 = _T_10366_number + _T_10368_number;
  assign _T_10396 = _T_10395[32:0];
  assign _T_10413 = _T_10364_number[7:0];
  assign _T_10415 = _T_10364_number[31:8];
  assign _T_10416 = {_T_10412,_T_10410};
  assign _T_10417 = x3437 ? x3455_number : x3450_number;
  assign _T_10418 = x3436 | x3437;
  assign _T_10433 = x3453_number[7:0];
  assign _T_10434 = x3453_number[31];
  assign _T_10435 = x3453_number[31:8];
  assign _T_10436 = {_T_10434,_T_10435};
  assign _T_10437 = {_T_10432,_T_10430};
  assign _T_10446 = x3456_number[7:0];
  assign _T_10447 = x3456_number[31];
  assign _T_10448 = x3456_number[31:8];
  assign _T_10449 = {_T_10447,_T_10448};
  assign _T_10450 = {_T_10445,_T_10443};
  assign _T_10451 = _T_10422_number + _T_10424_number;
  assign _T_10452 = _T_10451[32:0];
  assign _T_10469 = _T_10420_number[7:0];
  assign _T_10471 = _T_10420_number[31:8];
  assign _T_10472 = {_T_10468,_T_10466};
  assign _T_10473 = x3457 ? x3458_number : x3453_number;
  assign _T_10507 = _T_10482_number == 32'h0;
  assign _T_10522 = x3459_number[7:0];
  assign _T_10523 = x3459_number[31];
  assign _T_10524 = x3459_number[31:8];
  assign _T_10525 = {_T_10523,_T_10524};
  assign _T_10526 = {_T_10521,_T_10519};
  assign _T_10540 = _T_10511_number + 33'h0;
  assign _T_10541 = _T_10540[32:0];
  assign _T_10558 = _T_10509_number[7:0];
  assign _T_10560 = _T_10509_number[31:8];
  assign _T_10561 = {_T_10557,_T_10555};
  assign _T_10562 = x3462 ? x3459_number : x3463_number;
  assign _T_10565 = retime_released ? x3429_wren : 1'h0;
  assign _T_10568 = retime_released ? x3429_resetter : 1'h0;
  assign _T_10569 = reset | _T_10568;
  assign _T_10576 = retime_released ? _T_10574 : 1'h0;
  assign _T_10577 = b1204_chain_read_3 & _T_10576;
  assign _GEN_6 = {{2'd0}, x3305_number};
  assign _T_10600 = _GEN_6 << 2;
  assign x3308 = x3306_number[5:0];
  assign _GEN_7 = {{2'd0}, x3310_number};
  assign _T_10603 = _GEN_7 << 2;
  assign _T_10620 = x3306_number[31];
  assign _T_10622 = {_T_10620,x3306_number};
  assign _T_10633 = x3309_number[31];
  assign _T_10635 = {_T_10633,x3309_number};
  assign _T_10636 = _T_10607_number - _T_10609_number;
  assign _T_10637 = $unsigned(_T_10636);
  assign _T_10638 = _T_10637[32:0];
  assign _T_10658 = _T_10605_number[31:0];
  assign _T_10688 = x3311_number[31];
  assign _T_10690 = {_T_10688,x3311_number};
  assign _T_10691 = _T_10662_number + _T_10664_number;
  assign _T_10692 = _T_10691[32:0];
  assign _T_10712 = _T_10660_number[31:0];
  assign x3315 = x3313_number[5:0];
  assign _T_10743 = _T_10718_number == 32'h0;
  assign _T_10777 = x3316_number[31];
  assign _T_10779 = {_T_10777,x3316_number};
  assign _T_10780 = 33'h40 - _T_10753_number;
  assign _T_10781 = $unsigned(_T_10780);
  assign _T_10782 = _T_10781[32:0];
  assign _T_10802 = _T_10749_number[31:0];
  assign _T_10807 = x3317 ? 32'h0 : x3318_number;
  assign _T_10814 = _T_10633 ? 2'h3 : 2'h0;
  assign _T_10815 = x3309_number[31:2];
  assign _T_10816 = {_T_10814,_T_10815};
  assign _T_10819 = x3319_number[31];
  assign _T_10823 = _T_10819 ? 2'h3 : 2'h0;
  assign _T_10824 = x3319_number[31:2];
  assign _T_10825 = {_T_10823,_T_10824};
  assign _T_10842 = x3320_number[31];
  assign _T_10844 = {_T_10842,x3320_number};
  assign _T_10855 = x3310_number[31];
  assign _T_10857 = {_T_10855,x3310_number};
  assign _T_10858 = _T_10829_number + _T_10831_number;
  assign _T_10859 = _T_10858[32:0];
  assign _T_10879 = _T_10827_number[31:0];
  assign _T_10912 = _T_10883_number + _T_10885_number;
  assign _T_10913 = _T_10912[32:0];
  assign _T_10933 = _T_10881_number[31:0];
  assign _T_10950 = x3323_number[31];
  assign _T_10952 = {_T_10950,x3323_number};
  assign _T_10963 = x3321_number[31];
  assign _T_10965 = {_T_10963,x3321_number};
  assign _T_10966 = _T_10937_number + _T_10939_number;
  assign _T_10967 = _T_10966[32:0];
  assign _T_10987 = _T_10935_number[31:0];
  assign _T_11020 = _T_10991_number + _T_10993_number;
  assign _T_11021 = _T_11020[32:0];
  assign _T_11041 = _T_10989_number[31:0];
  assign _T_11058 = x3325_number[31];
  assign _T_11060 = {_T_11058,x3325_number};
  assign _T_11073 = {_T_10819,x3319_number};
  assign _T_11074 = _T_11045_number + _T_11047_number;
  assign _T_11075 = _T_11074[32:0];
  assign _T_11095 = _T_11043_number[31:0];
  assign _T_11106 = x3312_number[31];
  assign _T_11110 = _T_11106 ? 32'hffffffff : 32'h0;
  assign _T_11112 = {_T_11110,x3312_number};
  assign _T_11144 = x3327_number[63];
  assign _T_11146 = {_T_11144,x3327_number};
  assign _T_11157 = _T_11114_number[63];
  assign _T_11159 = {_T_11157,_T_11114_number};
  assign _T_11160 = _T_11131_number + _T_11133_number;
  assign _T_11161 = _T_11160[64:0];
  assign _T_11181 = _T_11129_number[63:0];
  assign _T_11194 = {1'h1,x3331_item1};
  assign _T_11195 = {_T_11194,x3331_item0};
  assign _T_11201 = retime_released ? x3335_datapath_en : 1'h0;
  assign _T_11202 = _T_11201 & b1204_chain_read_2;
  assign _T_11209 = b1204_chain_read_2 & _T_11201;
  assign _T_11210 = {x3333_item2,x3333_item1};
  assign _T_11211 = {_T_11210,x3333_item0};
  assign _T_11238 = retime_released ? x3283_datapath_en : 1'h0;
  assign _T_11239 = x3283_en & _T_11238;
  assign _T_11240 = _T_11239 & b1205_chain_read_1;
  assign _T_11254 = x3276[63:32];
  assign _T_11259 = b1205_chain_read_1 & _T_11238;
  assign _T_11264 = ~ _T_11259;
  assign _T_11265 = _T_11263 & _T_11264;
  assign _T_11266 = x3276[95:64];
  assign _T_11277 = _T_11275 & _T_11264;
  assign _T_11278 = x3276[31:0];
  assign _T_11289 = _T_11287 & _T_11264;
  assign _T_11306 = x3162_number[31];
  assign _T_11308 = {_T_11306,x3162_number};
  assign _T_11319 = b1202_number[31];
  assign _T_11321 = {_T_11319,b1202_number};
  assign _T_11322 = _T_11293_number - _T_11295_number;
  assign _T_11323 = $unsigned(_T_11322);
  assign _T_11324 = _T_11323[32:0];
  assign _T_11344 = _T_11291_number[31:0];
  assign _T_11376 = $signed(_T_11352_number);
  assign _T_11377 = $signed(32'sh40) < $signed(_T_11376);
  assign _T_11382_number = _T_11377 ? 32'h40 : x3163_number;
  assign _T_11440 = retime_released ? x3167_datapath_en : 1'h0;
  assign _T_11441 = b1204 & _T_11440;
  assign _T_11446 = ~ _T_11441;
  assign _T_11447 = _T_11445 & _T_11446;
  assign _T_11449 = x3410_en & retime_released;
  assign _T_11451 = x3410_sm_io_output_done;
  assign _T_11454 = x3410_sm_io_output_ctr_inc & _T_3809;
  assign _T_11455 = ~ x3410_ctr_trivial;
  assign _T_11456 = _T_11454 & _T_11455;
  assign _T_11457 = ~ x3410_sm_io_output_ctr_inc;
  assign _T_11466 = x3410_sm_io_output_ctr_inc & _T_11460;
  assign _T_11472 = retime_released ? _T_11470 : 1'h0;
  assign _T_11480 = retime_released ? _T_11478 : 1'h0;
  assign _T_11484 = $signed(x3411_number);
  assign _T_11753 = x3425_sm_io_output_done;
  assign _T_11755 = x3425_en & _T_3839;
  assign _T_11756 = ~ x3425_ctr_trivial;
  assign _T_11757 = _T_11755 & _T_11756;
  assign _T_11766 = retime_released ? _T_11764 : 1'h0;
  assign _T_11772 = retime_released ? _T_11770 : 1'h0;
  assign _T_11874 = $signed(_T_11849_number);
  assign _T_11875 = $signed(_T_11851_number);
  assign _T_11876 = $signed(_T_11874) < $signed(_T_11875);
  assign _T_11912 = retime_released ? _T_11910 : 1'h0;
  assign _T_11939 = _T_11914_number == 32'h0;
  assign _T_11940 = _T_11912 | _T_11939;
  assign _T_11941 = $unsigned(x3412_0);
  assign _T_11968 = $signed(_T_11943_number);
  assign _T_11969 = $signed(_T_11945_number);
  assign _T_11970 = $signed(_T_11968) <= $signed(_T_11969);
  assign _T_11997 = $signed(_T_11972_number);
  assign _T_11998 = $signed(_T_11974_number);
  assign _T_11999 = $signed(_T_11997) < $signed(_T_11998);
  assign _T_12000 = x3415 & x3417;
  assign _T_12017 = b1454_number[31];
  assign _T_12019 = {_T_12017,b1454_number};
  assign _T_12030 = x3414_number[31];
  assign _T_12032 = {_T_12030,x3414_number};
  assign _T_12033 = _T_12004_number - _T_12006_number;
  assign _T_12034 = $unsigned(_T_12033);
  assign _T_12035 = _T_12034[32:0];
  assign _T_12055 = _T_12002_number[31:0];
  assign _T_12056 = b1455 & b1205_chain_read_2;
  assign _T_12059 = x3420 & x3425_datapath_en;
  assign _T_12060 = x3418 & x3420;
  assign _T_12065 = x3423 & x3425_datapath_en;
  assign _T_12072 = retime_released ? x3220_datapath_en : 1'h0;
  assign _T_12073 = x3220_en & _T_12072;
  assign _T_12074 = _T_12073 & b1204_chain_read_1;
  assign _T_12088 = x3213[63:32];
  assign _T_12093 = b1204_chain_read_1 & _T_12072;
  assign _T_12098 = ~ _T_12093;
  assign _T_12099 = _T_12097 & _T_12098;
  assign _T_12100 = x3213[95:64];
  assign _T_12111 = _T_12109 & _T_12098;
  assign _T_12112 = x3213[31:0];
  assign _T_12123 = _T_12121 & _T_12098;
  assign _T_12124 = $unsigned(x3285_0);
  assign _T_12151 = $signed(_T_12126_number);
  assign _T_12152 = $signed(_T_12128_number);
  assign _T_12153 = $signed(_T_12151) <= $signed(_T_12152);
  assign _T_12180 = $signed(_T_12155_number);
  assign _T_12181 = $signed(_T_12157_number);
  assign _T_12182 = $signed(_T_12180) < $signed(_T_12181);
  assign _T_12183 = x3288 & x3290;
  assign _T_12200 = b1331_number[31];
  assign _T_12202 = {_T_12200,b1331_number};
  assign _T_12213 = x3287_number[31];
  assign _T_12215 = {_T_12213,x3287_number};
  assign _T_12216 = _T_12187_number - _T_12189_number;
  assign _T_12217 = $unsigned(_T_12216);
  assign _T_12218 = _T_12217[32:0];
  assign _T_12238 = _T_12185_number[31:0];
  assign _T_12239 = b1332 & b1205_chain_read_1;
  assign _T_12242 = x3293 & x3298_datapath_en;
  assign _T_12243 = x3291 & x3293;
  assign _T_12248 = x3296 & x3298_datapath_en;
  assign _T_12249 = $unsigned(x3222_0);
  assign _T_12276 = $signed(_T_12251_number);
  assign _T_12277 = $signed(_T_12253_number);
  assign _T_12278 = $signed(_T_12276) <= $signed(_T_12277);
  assign _T_12305 = $signed(_T_12280_number);
  assign _T_12306 = $signed(_T_12282_number);
  assign _T_12307 = $signed(_T_12305) < $signed(_T_12306);
  assign _T_12308 = x3225 & x3227;
  assign _T_12325 = b1270_number[31];
  assign _T_12327 = {_T_12325,b1270_number};
  assign _T_12338 = x3224_number[31];
  assign _T_12340 = {_T_12338,x3224_number};
  assign _T_12341 = _T_12312_number - _T_12314_number;
  assign _T_12342 = $unsigned(_T_12341);
  assign _T_12343 = _T_12342[32:0];
  assign _T_12363 = _T_12310_number[31:0];
  assign _T_12364 = b1271 & b1204_chain_read_1;
  assign _T_12367 = x3230 & x3235_datapath_en;
  assign _T_12368 = x3228 & x3230;
  assign _T_12373 = x3233 & x3235_datapath_en;
  assign _T_12380 = retime_released ? x3347_datapath_en : 1'h0;
  assign _T_12381 = x3347_en & _T_12380;
  assign _T_12382 = _T_12381 & b1204_chain_read_2;
  assign _T_12396 = x3340[63:32];
  assign _T_12401 = b1204_chain_read_2 & _T_12380;
  assign _T_12406 = ~ _T_12401;
  assign _T_12407 = _T_12405 & _T_12406;
  assign _T_12408 = x3340[95:64];
  assign _T_12419 = _T_12417 & _T_12406;
  assign _T_12420 = x3340[31:0];
  assign _T_12431 = _T_12429 & _T_12406;
  assign _T_12438 = retime_released ? x3410_datapath_en : 1'h0;
  assign _T_12439 = x3410_en & _T_12438;
  assign _T_12440 = _T_12439 & b1205_chain_read_2;
  assign _T_12454 = x3403[63:32];
  assign _T_12459 = b1205_chain_read_2 & _T_12438;
  assign _T_12464 = ~ _T_12459;
  assign _T_12465 = _T_12463 & _T_12464;
  assign _T_12466 = x3403[95:64];
  assign _T_12477 = _T_12475 & _T_12464;
  assign _T_12478 = x3403[31:0];
  assign _T_12489 = _T_12487 & _T_12464;
  assign io_done = done_latch_io_output_data;
  assign io_memStreams_loads_3_cmd_valid = x3365_valid;
  assign io_memStreams_loads_3_cmd_bits_addr = _T_3776;
  assign io_memStreams_loads_3_cmd_bits_isWr = _T_3779;
  assign io_memStreams_loads_3_cmd_bits_size = _T_3777[15:0];
  assign io_memStreams_loads_3_rdata_ready = x3367_ready;
  assign io_memStreams_loads_2_cmd_valid = x3302_valid;
  assign io_memStreams_loads_2_cmd_bits_addr = _T_9360;
  assign io_memStreams_loads_2_cmd_bits_isWr = _T_9363;
  assign io_memStreams_loads_2_cmd_bits_size = _T_9361[15:0];
  assign io_memStreams_loads_2_rdata_ready = x3304_ready;
  assign io_memStreams_loads_1_cmd_valid = x3238_valid;
  assign io_memStreams_loads_1_cmd_bits_addr = _T_4545;
  assign io_memStreams_loads_1_cmd_bits_isWr = _T_4548;
  assign io_memStreams_loads_1_cmd_bits_size = _T_4546[15:0];
  assign io_memStreams_loads_1_rdata_ready = x3240_ready;
  assign io_memStreams_loads_0_cmd_valid = x3175_valid;
  assign io_memStreams_loads_0_cmd_bits_addr = _T_3026;
  assign io_memStreams_loads_0_cmd_bits_isWr = _T_3029;
  assign io_memStreams_loads_0_cmd_bits_size = _T_3027[15:0];
  assign io_memStreams_loads_0_rdata_ready = x3177_ready;
  assign io_argOuts_0_valid = x3141_en_options_0;
  assign io_argOuts_0_bits = x3141_data_options_0;
  assign x3141_data_options_0 = _T_7015;
  assign x3141_en_options_0 = x3518_datapath_en;
  assign RootController_done = _T_1688;
  assign RootController_en = _T_1698;
  assign RootController_resetter = _T_1702;
  assign RetimeWrapper_io_flow = 1'h1;
  assign RetimeWrapper_io_in = 1'h0;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign retime_released = _T_1710;
  assign x3153_number = io_argIns_0[31:0];
  assign x3155_en = _T_1996;
  assign x3155_resetter = _T_1999;
  assign x3154_0 = x3155_io_output_counts_0;
  assign x3154_1 = x3155_io_output_counts_1;
  assign x3515_level0_iters = _T_1964_number;
  assign x3515_done = _T_1991;
  assign x3515_en = x3515_base_en;
  assign x3515_base_en = _T_2486;
  assign x3515_resetter = _T_2492;
  assign x3515_ctr_trivial = _T_2424;
  assign x3515_rst_en = x3515_sm_io_output_rst_en;
  assign x3152_wren = x3514_sm_io_output_done;
  assign x3152_resetter = x3515_rst_en;
  assign b1202_number = _T_2513;
  assign b1203_number = _T_2514;
  assign x3174_done = _T_2530;
  assign x3174_en = x3174_base_en;
  assign x3174_base_en = _T_2290;
  assign x3174_resetter = _T_2296;
  assign x3174_ctr_trivial = _T_2543;
  assign x3167_done = _T_8330;
  assign x3167_en = x3167_base_en;
  assign x3167_base_en = _T_2559;
  assign x3167_mask = b1204;
  assign x3167_resetter = _T_2565;
  assign x3167_datapath_en = _T_8335;
  assign x3167_ctr_trivial = _T_8359;
  assign x3162_number = io_argIns_0[31:0];
  assign x3163_number = _T_11326_number;
  assign x3164_number = _T_11382_number;
  assign x3173_done = _T_8376;
  assign x3173_en = x3173_base_en;
  assign x3173_base_en = _T_2579;
  assign x3173_mask = b1205;
  assign x3173_resetter = _T_2585;
  assign x3173_datapath_en = _T_8381;
  assign x3173_ctr_trivial = _T_8405;
  assign x3168_number = io_argIns_0[31:0];
  assign x3169_number = _T_8445_number;
  assign x3170_number = _T_8501_number;
  assign x3301_done = _T_2600;
  assign x3301_en = x3301_base_en;
  assign x3301_base_en = _T_2310;
  assign x3301_resetter = _T_2316;
  assign x3301_ctr_trivial = _T_2613;
  assign x3237_done = _T_2848;
  assign x3237_en = x3237_base_en;
  assign x3237_base_en = _T_2629;
  assign x3237_mask = b1204_chain_read_1;
  assign x3237_resetter = _T_2635;
  assign x3237_ctr_trivial = _T_2861;
  assign x3175_valid_options_0 = _T_4473;
  assign x3175_valid_stops_0 = x3208_done;
  assign x3175_valid = _T_4480;
  assign x3175_data_options_0 = x3204;
  assign x3175_ready = _T_3025;
  assign x3177_ready_options_0 = _T_12367;
  assign x3177_ready = x3177_ready_options_0;
  assign x3177_now_valid = io_memStreams_loads_0_rdata_valid;
  assign x3177_valid = _T_3034;
  assign x3177_0_number = io_memStreams_loads_0_rdata_bits_0;
  assign x3208_done = _T_2987;
  assign x3208_en = _T_2888;
  assign x3208_base_en = _T_2877;
  assign x3208_mask = b1204_chain_read_1;
  assign x3208_resetter = _T_2894;
  assign x3208_datapath_en = _T_2992;
  assign x3208_ctr_trivial = _T_3018;
  assign x3178_number = _T_3855_number;
  assign x3179_number = _T_3870_number;
  assign x3182_number = {{26'd0}, x3181};
  assign x3183_number = x3156_0_io_output_1_data;
  assign x3184_number = _T_3873_number;
  assign x3185_number = _T_3911_number;
  assign x3186_number = _T_3965_number;
  assign x3189_number = {{26'd0}, x3188};
  assign x3190 = _T_4014;
  assign x3191_number = _T_4055_number;
  assign x3192_number = _T_4078;
  assign x3193_number = _T_4080_number;
  assign x3194_number = _T_4089_number;
  assign x3195_number = _T_4132_number;
  assign x3196_number = _T_4186_number;
  assign x3197_number = _T_4240_number;
  assign x3198_number = _T_4294_number;
  assign x3199_number = _T_4348_number;
  assign x3200_number = _T_4374;
  assign x3202_number = _T_4434_number;
  assign x3203_number = _T_4460;
  assign x3204_item0 = x3203_number;
  assign x3204_item1 = x3199_number;
  assign x3204 = _T_4466;
  assign x3206_item0 = x3197_number;
  assign x3206_item1 = x3193_number;
  assign x3206_item2 = x3195_number;
  assign x3206 = _T_4482;
  assign x3236_done = _T_3037;
  assign x3236_en = x3236_base_en;
  assign x3236_base_en = _T_2908;
  assign x3236_mask = b1204_chain_read_1;
  assign x3236_resetter = _T_2914;
  assign x3236_ctr_trivial = _T_3050;
  assign x3220_done = _T_3106;
  assign x3220_en = _T_3076;
  assign x3220_base_en = _T_3066;
  assign x3220_mask = b1204_chain_read_1;
  assign x3220_resetter = _T_3082;
  assign x3220_datapath_en = _T_3111;
  assign x3220_ctr_trivial = _T_3135;
  assign x3214_number = _T_12088;
  assign x3216_number = _T_12100;
  assign x3218_number = _T_12112;
  assign x3221_number = x3212_0_io_output_data;
  assign x3223_done = x3223_io_output_done;
  assign x3223_en = x3235_datapath_en;
  assign x3223_resetter = _T_3421;
  assign x3222_0 = x3223_io_output_counts_0;
  assign x3235_done = _T_3408;
  assign x3235_en = _T_3097;
  assign x3235_base_en = _T_3096;
  assign x3235_mask = b1204_chain_read_1;
  assign x3235_datapath_en = _T_3412;
  assign x3235_ctr_trivial = _T_3595;
  assign b1270_number = _T_12249;
  assign x3224_number = x3210_0_io_output_data;
  assign x3225 = _T_12278;
  assign x3226_number = x3211_0_io_output_data;
  assign x3227 = _T_12307;
  assign x3228 = _T_12308;
  assign x3229_number = _T_12345_number;
  assign x3230 = _T_12364;
  assign x3232_number = x3177_0_number;
  assign x3233 = _T_12368;
  assign x3234_wVec_0_addr_0 = x3229_number[5:0];
  assign x3234_wVec_0_data = x3232_number;
  assign x3234_wVec_0_en = _T_12373;
  assign x3300_done = _T_2917;
  assign x3300_en = x3300_base_en;
  assign x3300_base_en = _T_2649;
  assign x3300_mask = b1205_chain_read_1;
  assign x3300_resetter = _T_2655;
  assign x3300_ctr_trivial = _T_2930;
  assign x3238_valid_options_0 = _T_7638;
  assign x3238_valid_stops_0 = x3271_done;
  assign x3238_valid = _T_7645;
  assign x3238_data_options_0 = x3267;
  assign x3238_ready = _T_4544;
  assign x3240_ready_options_0 = _T_12242;
  assign x3240_ready = x3240_ready_options_0;
  assign x3240_now_valid = io_memStreams_loads_1_rdata_valid;
  assign x3240_valid = _T_4553;
  assign x3240_0_number = io_memStreams_loads_1_rdata_bits_0;
  assign x3271_done = _T_4506;
  assign x3271_en = _T_2957;
  assign x3271_base_en = _T_2946;
  assign x3271_mask = b1205_chain_read_1;
  assign x3271_resetter = _T_2963;
  assign x3271_datapath_en = _T_4511;
  assign x3271_ctr_trivial = _T_4537;
  assign x3241_number = _T_7020_number;
  assign x3242_number = _T_7035_number;
  assign x3245_number = {{26'd0}, x3244};
  assign x3246_number = x3157_0_io_output_1_data;
  assign x3247_number = _T_7038_number;
  assign x3248_number = _T_7076_number;
  assign x3249_number = _T_7130_number;
  assign x3252_number = {{26'd0}, x3251};
  assign x3253 = _T_7179;
  assign x3254_number = _T_7220_number;
  assign x3255_number = _T_7243;
  assign x3256_number = _T_7245_number;
  assign x3257_number = _T_7254_number;
  assign x3258_number = _T_7297_number;
  assign x3259_number = _T_7351_number;
  assign x3260_number = _T_7405_number;
  assign x3261_number = _T_7459_number;
  assign x3262_number = _T_7513_number;
  assign x3263_number = _T_7539;
  assign x3265_number = _T_7599_number;
  assign x3266_number = _T_7625;
  assign x3267_item0 = x3266_number;
  assign x3267_item1 = x3262_number;
  assign x3267 = _T_7631;
  assign x3269_item0 = x3260_number;
  assign x3269_item1 = x3256_number;
  assign x3269_item2 = x3258_number;
  assign x3269 = _T_7647;
  assign x3299_done = _T_4556;
  assign x3299_en = x3299_base_en;
  assign x3299_base_en = _T_2977;
  assign x3299_mask = b1205_chain_read_1;
  assign x3299_resetter = _T_2983;
  assign x3299_ctr_trivial = _T_4569;
  assign x3283_done = _T_4625;
  assign x3283_en = _T_4595;
  assign x3283_base_en = _T_4585;
  assign x3283_mask = b1205_chain_read_1;
  assign x3283_resetter = _T_4601;
  assign x3283_datapath_en = _T_4630;
  assign x3283_ctr_trivial = _T_4654;
  assign x3277_number = _T_11254;
  assign x3279_number = _T_11266;
  assign x3281_number = _T_11278;
  assign x3284_number = x3275_0_io_output_data;
  assign x3286_done = x3286_io_output_done;
  assign x3286_en = x3298_datapath_en;
  assign x3286_resetter = _T_4940;
  assign x3285_0 = x3286_io_output_counts_0;
  assign x3298_done = _T_4927;
  assign x3298_en = _T_4616;
  assign x3298_base_en = _T_4615;
  assign x3298_mask = b1205_chain_read_1;
  assign x3298_datapath_en = _T_4931;
  assign x3298_ctr_trivial = _T_5114;
  assign b1331_number = _T_12124;
  assign x3287_number = x3273_0_io_output_data;
  assign x3288 = _T_12153;
  assign x3289_number = x3274_0_io_output_data;
  assign x3290 = _T_12182;
  assign x3291 = _T_12183;
  assign x3292_number = _T_12220_number;
  assign x3293 = _T_12239;
  assign x3295_number = x3240_0_number;
  assign x3296 = _T_12243;
  assign x3297_wVec_0_addr_0 = x3292_number[5:0];
  assign x3297_wVec_0_data = x3295_number;
  assign x3297_wVec_0_en = _T_12248;
  assign x3428_done = _T_2670;
  assign x3428_en = x3428_base_en;
  assign x3428_base_en = _T_2330;
  assign x3428_resetter = _T_2336;
  assign x3428_ctr_trivial = _T_2683;
  assign x3364_done = _T_3598;
  assign x3364_en = x3364_base_en;
  assign x3364_base_en = _T_2699;
  assign x3364_mask = b1204_chain_read_2;
  assign x3364_resetter = _T_2705;
  assign x3364_ctr_trivial = _T_3611;
  assign x3302_valid_options_0 = _T_11202;
  assign x3302_valid_stops_0 = x3335_done;
  assign x3302_valid = _T_11209;
  assign x3302_data_options_0 = x3331;
  assign x3302_ready = _T_9359;
  assign x3304_ready_options_0 = _T_10048;
  assign x3304_ready = x3304_ready_options_0;
  assign x3304_now_valid = io_memStreams_loads_2_rdata_valid;
  assign x3304_valid = _T_9368;
  assign x3304_0_number = io_memStreams_loads_2_rdata_bits_0;
  assign x3335_done = _T_9321;
  assign x3335_en = _T_3638;
  assign x3335_base_en = _T_3627;
  assign x3335_mask = b1204_chain_read_2;
  assign x3335_resetter = _T_3644;
  assign x3335_datapath_en = _T_9326;
  assign x3335_ctr_trivial = _T_9352;
  assign x3305_number = _T_10584_number;
  assign x3306_number = _T_10599_number;
  assign x3309_number = {{26'd0}, x3308};
  assign x3310_number = x3156_0_io_output_2_data;
  assign x3311_number = _T_10602_number;
  assign x3312_number = _T_10640_number;
  assign x3313_number = _T_10694_number;
  assign x3316_number = {{26'd0}, x3315};
  assign x3317 = _T_10743;
  assign x3318_number = _T_10784_number;
  assign x3319_number = _T_10807;
  assign x3320_number = _T_10809_number;
  assign x3321_number = _T_10818_number;
  assign x3322_number = _T_10861_number;
  assign x3323_number = _T_10915_number;
  assign x3324_number = _T_10969_number;
  assign x3325_number = _T_11023_number;
  assign x3326_number = _T_11077_number;
  assign x3327_number = _T_11103;
  assign x3329_number = _T_11163_number;
  assign x3330_number = _T_11189;
  assign x3331_item0 = x3330_number;
  assign x3331_item1 = x3326_number;
  assign x3331 = _T_11195;
  assign x3333_item0 = x3324_number;
  assign x3333_item1 = x3320_number;
  assign x3333_item2 = x3322_number;
  assign x3333 = _T_11211;
  assign x3363_done = _T_9371;
  assign x3363_en = x3363_base_en;
  assign x3363_base_en = _T_3658;
  assign x3363_mask = b1204_chain_read_2;
  assign x3363_resetter = _T_3664;
  assign x3363_ctr_trivial = _T_9384;
  assign x3347_done = _T_9440;
  assign x3347_en = _T_9410;
  assign x3347_base_en = _T_9400;
  assign x3347_mask = b1204_chain_read_2;
  assign x3347_resetter = _T_9416;
  assign x3347_datapath_en = _T_9445;
  assign x3347_ctr_trivial = _T_9469;
  assign x3341_number = _T_12396;
  assign x3343_number = _T_12408;
  assign x3345_number = _T_12420;
  assign x3348_number = x3339_0_io_output_data;
  assign x3350_done = x3350_io_output_done;
  assign x3350_en = x3362_datapath_en;
  assign x3350_resetter = _T_9755;
  assign x3349_0 = x3350_io_output_counts_0;
  assign x3362_done = _T_9742;
  assign x3362_en = _T_9431;
  assign x3362_base_en = _T_9430;
  assign x3362_mask = b1204_chain_read_2;
  assign x3362_datapath_en = _T_9746;
  assign x3362_ctr_trivial = _T_9929;
  assign b1393_number = _T_9930;
  assign x3351_number = x3337_0_io_output_data;
  assign x3352 = _T_9959;
  assign x3353_number = x3338_0_io_output_data;
  assign x3354 = _T_9988;
  assign x3355 = _T_9989;
  assign x3356_number = _T_10026_number;
  assign x3357 = _T_10045;
  assign x3359_number = x3304_0_number;
  assign x3360 = _T_10049;
  assign x3361_wVec_0_addr_0 = x3356_number[5:0];
  assign x3361_wVec_0_data = x3359_number;
  assign x3361_wVec_0_en = _T_10054;
  assign x3427_done = _T_3667;
  assign x3427_en = x3427_base_en;
  assign x3427_base_en = _T_2719;
  assign x3427_mask = b1205_chain_read_2;
  assign x3427_resetter = _T_2725;
  assign x3427_ctr_trivial = _T_3680;
  assign x3365_valid_options_0 = _T_8287;
  assign x3365_valid_stops_0 = x3398_done;
  assign x3365_valid = _T_8294;
  assign x3365_data_options_0 = x3394;
  assign x3365_ready = _T_3775;
  assign x3367_ready_options_0 = _T_12059;
  assign x3367_ready = x3367_ready_options_0;
  assign x3367_now_valid = io_memStreams_loads_3_rdata_valid;
  assign x3367_valid = _T_3784;
  assign x3367_0_number = io_memStreams_loads_3_rdata_bits_0;
  assign x3398_done = _T_3737;
  assign x3398_en = _T_3707;
  assign x3398_base_en = _T_3696;
  assign x3398_mask = b1205_chain_read_2;
  assign x3398_resetter = _T_3713;
  assign x3398_datapath_en = _T_3742;
  assign x3398_ctr_trivial = _T_3768;
  assign x3368_number = _T_7669_number;
  assign x3369_number = _T_7684_number;
  assign x3372_number = {{26'd0}, x3371};
  assign x3373_number = x3157_0_io_output_2_data;
  assign x3374_number = _T_7687_number;
  assign x3375_number = _T_7725_number;
  assign x3376_number = _T_7779_number;
  assign x3379_number = {{26'd0}, x3378};
  assign x3380 = _T_7828;
  assign x3381_number = _T_7869_number;
  assign x3382_number = _T_7892;
  assign x3383_number = _T_7894_number;
  assign x3384_number = _T_7903_number;
  assign x3385_number = _T_7946_number;
  assign x3386_number = _T_8000_number;
  assign x3387_number = _T_8054_number;
  assign x3388_number = _T_8108_number;
  assign x3389_number = _T_8162_number;
  assign x3390_number = _T_8188;
  assign x3392_number = _T_8248_number;
  assign x3393_number = _T_8274;
  assign x3394_item0 = x3393_number;
  assign x3394_item1 = x3389_number;
  assign x3394 = _T_8280;
  assign x3396_item0 = x3387_number;
  assign x3396_item1 = x3383_number;
  assign x3396_item2 = x3385_number;
  assign x3396 = _T_8296;
  assign x3426_done = _T_3787;
  assign x3426_en = x3426_base_en;
  assign x3426_base_en = _T_3727;
  assign x3426_mask = b1205_chain_read_2;
  assign x3426_resetter = _T_3733;
  assign x3426_ctr_trivial = _T_3800;
  assign x3410_done = _T_11451;
  assign x3410_en = _T_3826;
  assign x3410_base_en = _T_3816;
  assign x3410_mask = b1205_chain_read_2;
  assign x3410_resetter = _T_3832;
  assign x3410_datapath_en = _T_11456;
  assign x3410_ctr_trivial = _T_11480;
  assign x3404_number = _T_12454;
  assign x3406_number = _T_12466;
  assign x3408_number = _T_12478;
  assign x3411_number = x3402_0_io_output_data;
  assign x3413_done = x3413_io_output_done;
  assign x3413_en = x3425_datapath_en;
  assign x3413_resetter = _T_11766;
  assign x3412_0 = x3413_io_output_counts_0;
  assign x3425_done = _T_11753;
  assign x3425_en = _T_3847;
  assign x3425_base_en = _T_3846;
  assign x3425_mask = b1205_chain_read_2;
  assign x3425_datapath_en = _T_11757;
  assign x3425_ctr_trivial = _T_11940;
  assign b1454_number = _T_11941;
  assign x3414_number = x3400_0_io_output_data;
  assign x3415 = _T_11970;
  assign x3416_number = x3401_0_io_output_data;
  assign x3417 = _T_11999;
  assign x3418 = _T_12000;
  assign x3419_number = _T_12037_number;
  assign x3420 = _T_12056;
  assign x3422_number = x3367_0_number;
  assign x3423 = _T_12060;
  assign x3424_wVec_0_addr_0 = x3419_number[5:0];
  assign x3424_wVec_0_data = x3422_number;
  assign x3424_wVec_0_en = _T_12065;
  assign x3503_done = _T_2742;
  assign x3503_en = x3503_base_en;
  assign x3503_base_en = _T_2350;
  assign x3503_resetter = _T_2356;
  assign x3503_ctr_trivial = _T_2755;
  assign x3431_number = x3156_0_io_output_3_data;
  assign x3433_done = x3433_io_output_done;
  assign x3433_en = _T_5400;
  assign x3433_resetter = _T_5403;
  assign x3432_0 = x3433_io_output_counts_0;
  assign x3432_1 = x3433_io_output_counts_1;
  assign x3432_2 = x3433_io_output_counts_2;
  assign x3432_3 = x3433_io_output_counts_3;
  assign x3466_done = _T_5395;
  assign x3466_en = x3466_base_en;
  assign x3466_base_en = _T_2771;
  assign x3466_mask = b1204_chain_read_3;
  assign x3466_resetter = _T_2777;
  assign x3466_datapath_en = _T_5399;
  assign x3466_ctr_trivial = _T_5972;
  assign x3466_rst_en = x3466_sm_io_output_rst_en;
  assign x3429_wren = _T_5416;
  assign x3429_resetter = x3466_rst_en;
  assign b1479_number = _T_10055;
  assign b1480_number = _T_10056;
  assign b1481_number = _T_10057;
  assign b1482_number = _T_10058;
  assign x3434 = _T_10059;
  assign x3435 = _T_10060;
  assign x3436 = _T_10061;
  assign x3437 = _T_10062;
  assign x3438_rVec_0_addr_0 = b1479_number[5:0];
  assign x3438_rVec_0_en = _T_10066;
  assign x3438_rVec_1_addr_0 = b1480_number[5:0];
  assign x3438_rVec_1_en = _T_10070;
  assign x3438_rVec_2_addr_0 = b1481_number[5:0];
  assign x3438_rVec_2_en = _T_10074;
  assign x3438_rVec_3_addr_0 = b1482_number[5:0];
  assign x3438_rVec_3_en = _T_10078;
  assign x3439_number = x3438_0_number;
  assign x3440_number = x3438_1_number;
  assign x3441_number = x3438_2_number;
  assign x3442_number = x3438_3_number;
  assign x3443_rVec_0_addr_0 = b1479_number[5:0];
  assign x3443_rVec_0_en = _T_10066;
  assign x3443_rVec_1_addr_0 = b1480_number[5:0];
  assign x3443_rVec_1_en = _T_10070;
  assign x3443_rVec_2_addr_0 = b1481_number[5:0];
  assign x3443_rVec_2_en = _T_10074;
  assign x3443_rVec_3_addr_0 = b1482_number[5:0];
  assign x3443_rVec_3_en = _T_10078;
  assign x3444_number = x3443_0_number;
  assign x3445_number = x3443_1_number;
  assign x3446_number = x3443_2_number;
  assign x3447_number = x3443_3_number;
  assign x3448_number = _T_10180_number;
  assign x3449_number = _T_10216_number;
  assign x3450_number = _T_10252_number;
  assign x3451_number = _T_10288_number;
  assign x3452_number = _T_10342_number;
  assign x3453_number = _T_10361;
  assign x3455_number = _T_10398_number;
  assign x3456_number = _T_10417;
  assign x3457 = _T_10418;
  assign x3458_number = _T_10454_number;
  assign x3459_number = _T_10473;
  assign x3462 = _T_10507;
  assign x3463_number = _T_10543_number;
  assign x3464_number = _T_10562;
  assign x3465_number = x3429_0_io_output;
  assign x3467_number = x3157_0_io_output_3_data;
  assign x3469_done = x3469_io_output_done;
  assign x3469_en = _T_6258;
  assign x3469_resetter = _T_6261;
  assign x3468_0 = x3469_io_output_counts_0;
  assign x3468_1 = x3469_io_output_counts_1;
  assign x3468_2 = x3469_io_output_counts_2;
  assign x3468_3 = x3469_io_output_counts_3;
  assign x3502_done = _T_6253;
  assign x3502_en = x3502_base_en;
  assign x3502_base_en = _T_2791;
  assign x3502_mask = b1205_chain_read_3;
  assign x3502_resetter = _T_2797;
  assign x3502_datapath_en = _T_6257;
  assign x3502_ctr_trivial = _T_6830;
  assign x3502_rst_en = x3502_sm_io_output_rst_en;
  assign x3430_wren = _T_6274;
  assign x3430_resetter = x3502_rst_en;
  assign b1520_number = _T_8790;
  assign b1521_number = _T_8791;
  assign b1522_number = _T_8792;
  assign b1523_number = _T_8793;
  assign x3470 = _T_8794;
  assign x3471 = _T_8795;
  assign x3472 = _T_8796;
  assign x3473 = _T_8797;
  assign x3474_rVec_0_addr_0 = b1520_number[5:0];
  assign x3474_rVec_0_en = _T_8801;
  assign x3474_rVec_1_addr_0 = b1521_number[5:0];
  assign x3474_rVec_1_en = _T_8805;
  assign x3474_rVec_2_addr_0 = b1522_number[5:0];
  assign x3474_rVec_2_en = _T_8809;
  assign x3474_rVec_3_addr_0 = b1523_number[5:0];
  assign x3474_rVec_3_en = _T_8813;
  assign x3475_number = x3474_0_number;
  assign x3476_number = x3474_1_number;
  assign x3477_number = x3474_2_number;
  assign x3478_number = x3474_3_number;
  assign x3479_rVec_0_addr_0 = b1520_number[5:0];
  assign x3479_rVec_0_en = _T_8801;
  assign x3479_rVec_1_addr_0 = b1521_number[5:0];
  assign x3479_rVec_1_en = _T_8805;
  assign x3479_rVec_2_addr_0 = b1522_number[5:0];
  assign x3479_rVec_2_en = _T_8809;
  assign x3479_rVec_3_addr_0 = b1523_number[5:0];
  assign x3479_rVec_3_en = _T_8813;
  assign x3480_number = x3479_0_number;
  assign x3481_number = x3479_1_number;
  assign x3482_number = x3479_2_number;
  assign x3483_number = x3479_3_number;
  assign x3484_number = _T_8915_number;
  assign x3485_number = _T_8951_number;
  assign x3486_number = _T_8987_number;
  assign x3487_number = _T_9023_number;
  assign x3488_number = _T_9077_number;
  assign x3489_number = _T_9096;
  assign x3491_number = _T_9133_number;
  assign x3492_number = _T_9152;
  assign x3493 = _T_9153;
  assign x3494_number = _T_9189_number;
  assign x3495_number = _T_9208;
  assign x3498 = _T_9242;
  assign x3499_number = _T_9278_number;
  assign x3500_number = _T_9297;
  assign x3501_number = x3430_0_io_output;
  assign x3514_done = _T_2812;
  assign x3514_en = x3514_base_en;
  assign x3514_base_en = _T_2370;
  assign x3514_resetter = _T_2376;
  assign x3504_number = x3430_1_io_output_1_data;
  assign x3505_number = x3429_1_io_output_1_data;
  assign x3506_number = _T_6866_number;
  assign x3507_number = _T_6885;
  assign x3510 = _T_6934;
  assign x3511_number = _T_6970_number;
  assign x3512_number = _T_6989;
  assign x3513_number = x3152_1_io_output;
  assign x3518_done = _T_2439;
  assign x3518_en = x3518_base_en;
  assign x3518_base_en = _T_2506;
  assign x3518_resetter = _T_2512;
  assign x3518_datapath_en = _T_2444;
  assign x3518_ctr_trivial = _T_2468;
  assign x3516_number = x3152_0_io_output_data;
  assign RootController_sm_io_input_enable = _T_1675;
  assign RootController_sm_io_input_stageDone_0 = x3515_done;
  assign RootController_sm_io_input_stageDone_1 = x3518_done;
  assign RootController_sm_io_input_stageMask_0 = 1'h1;
  assign RootController_sm_io_input_stageMask_1 = 1'h1;
  assign RootController_sm_io_input_rst = RootController_resetter;
  assign RootController_sm_clock = clock;
  assign RootController_sm_reset = reset;
  assign x3152_0_io_input_0_data = x3513_number;
  assign x3152_0_io_input_0_init = 32'h0;
  assign x3152_0_io_input_0_enable = _T_6997;
  assign x3152_0_io_input_0_reset = _T_7002;
  assign x3152_0_clock = clock;
  assign x3152_0_reset = reset;
  assign x3152_1_io_input_next = x3512_number;
  assign x3152_1_io_input_enable = _T_7005;
  assign x3152_1_io_input_reset = _T_7009;
  assign x3152_1_clock = clock;
  assign x3152_1_reset = reset;
  assign x3155_io_input_stops_0 = _T_1711;
  assign x3155_io_input_reset = x3155_resetter;
  assign x3155_io_input_enable = x3155_en;
  assign x3155_clock = clock;
  assign x3155_reset = reset;
  assign x3515_sm_io_input_enable = _T_1978;
  assign x3515_sm_io_input_numIter = x3515_level0_iters;
  assign x3515_sm_io_input_stageDone_0 = x3174_done;
  assign x3515_sm_io_input_stageDone_1 = x3301_done;
  assign x3515_sm_io_input_stageDone_2 = x3428_done;
  assign x3515_sm_io_input_stageDone_3 = x3503_done;
  assign x3515_sm_io_input_stageDone_4 = x3514_done;
  assign x3515_sm_io_input_rst = x3515_resetter;
  assign x3515_sm_clock = clock;
  assign x3515_sm_reset = reset;
  assign b1204 = _T_2102;
  assign b1204_chain_read_1 = _T_1660;
  assign b1204_chain_read_2 = _T_1662;
  assign b1204_chain_read_3 = _T_1664;
  assign b1205 = _T_2239;
  assign b1205_chain_read_1 = _T_1668;
  assign b1205_chain_read_2 = _T_1670;
  assign b1205_chain_read_3 = _T_1672;
  assign b1205_chain_read_4 = _T_1674;
  assign b1202_chain_io_sEn_0 = x3174_en;
  assign b1202_chain_io_sEn_1 = x3301_en;
  assign b1202_chain_io_sEn_2 = x3428_en;
  assign b1202_chain_io_sEn_3 = x3503_en;
  assign b1202_chain_io_sEn_4 = x3514_en;
  assign b1202_chain_io_sDone_0 = _T_8630;
  assign b1202_chain_io_sDone_1 = _T_8633;
  assign b1202_chain_io_sDone_2 = _T_8636;
  assign b1202_chain_io_sDone_3 = _T_8639;
  assign b1202_chain_io_sDone_4 = _T_8642;
  assign b1202_chain_io_input_0_data = b1202_number;
  assign b1202_chain_io_input_0_enable = x3515_sm_io_output_ctr_inc;
  assign b1202_chain_io_input_0_reset = _T_2380;
  assign b1202_chain_clock = clock;
  assign b1202_chain_reset = reset;
  assign b1202_chain_read_1 = b1202_chain_io_output_1_data;
  assign b1202_chain_read_2 = b1202_chain_io_output_2_data;
  assign b1202_chain_read_4 = b1202_chain_io_output_4_data;
  assign b1203_chain_io_sEn_0 = x3174_en;
  assign b1203_chain_io_sEn_1 = x3301_en;
  assign b1203_chain_io_sEn_2 = x3428_en;
  assign b1203_chain_io_sEn_3 = x3503_en;
  assign b1203_chain_io_sEn_4 = x3514_en;
  assign b1203_chain_io_sDone_0 = _T_8630;
  assign b1203_chain_io_sDone_1 = _T_8633;
  assign b1203_chain_io_sDone_2 = _T_8636;
  assign b1203_chain_io_sDone_3 = _T_8639;
  assign b1203_chain_io_sDone_4 = _T_8642;
  assign b1203_chain_io_input_0_data = b1203_number;
  assign b1203_chain_io_input_0_enable = x3515_sm_io_output_ctr_inc;
  assign b1203_chain_io_input_0_reset = _T_2387;
  assign b1203_chain_clock = clock;
  assign b1203_chain_reset = reset;
  assign b1203_chain_read_1 = b1203_chain_io_output_1_data;
  assign b1203_chain_read_2 = b1203_chain_io_output_2_data;
  assign x3156_0_io_sEn_0 = x3174_base_en;
  assign x3156_0_io_sEn_1 = x3301_base_en;
  assign x3156_0_io_sEn_2 = x3428_base_en;
  assign x3156_0_io_sEn_3 = x3503_base_en;
  assign x3156_0_io_sDone_0 = _T_8663;
  assign x3156_0_io_sDone_1 = _T_8669;
  assign x3156_0_io_sDone_2 = _T_8675;
  assign x3156_0_io_sDone_3 = _T_8681;
  assign x3156_0_io_input_0_data = x3164_number;
  assign x3156_0_io_input_0_enable = _T_11441;
  assign x3156_0_io_input_0_reset = _T_11447;
  assign x3156_0_clock = clock;
  assign x3156_0_reset = reset;
  assign x3157_0_io_sEn_0 = x3174_base_en;
  assign x3157_0_io_sEn_1 = x3301_base_en;
  assign x3157_0_io_sEn_2 = x3428_base_en;
  assign x3157_0_io_sEn_3 = x3503_base_en;
  assign x3157_0_io_sDone_0 = _T_8687;
  assign x3157_0_io_sDone_1 = _T_8693;
  assign x3157_0_io_sDone_2 = _T_8699;
  assign x3157_0_io_sDone_3 = _T_8705;
  assign x3157_0_io_input_0_data = x3170_number;
  assign x3157_0_io_input_0_enable = _T_8560;
  assign x3157_0_io_input_0_reset = _T_8566;
  assign x3157_0_clock = clock;
  assign x3157_0_reset = reset;
  assign x3158_0_io_sEn_0 = x3301_base_en;
  assign x3158_0_io_sEn_1 = x3428_base_en;
  assign x3158_0_io_sEn_2 = x3503_base_en;
  assign x3158_0_io_sDone_0 = _T_8735;
  assign x3158_0_io_sDone_1 = _T_8741;
  assign x3158_0_io_sDone_2 = _T_8747;
  assign x3158_0_io_w_0_addr_0 = x3234_wVec_0_addr_0;
  assign x3158_0_io_w_0_data = x3234_wVec_0_data;
  assign x3158_0_io_w_0_en = x3234_wVec_0_en;
  assign x3158_0_io_r_0_addr_0 = _T_10086_0_addr_0;
  assign x3158_0_io_r_0_en = _T_10086_0_en;
  assign x3158_0_io_r_1_addr_0 = _T_10086_1_addr_0;
  assign x3158_0_io_r_1_en = _T_10086_1_en;
  assign x3158_0_io_r_2_addr_0 = _T_10086_2_addr_0;
  assign x3158_0_io_r_2_en = _T_10086_2_en;
  assign x3158_0_io_r_3_addr_0 = _T_10086_3_addr_0;
  assign x3158_0_io_r_3_en = _T_10086_3_en;
  assign x3158_0_clock = clock;
  assign x3158_0_reset = reset;
  assign x3159_0_io_sEn_0 = x3301_base_en;
  assign x3159_0_io_sEn_1 = x3428_base_en;
  assign x3159_0_io_sEn_2 = x3503_base_en;
  assign x3159_0_io_sDone_0 = _T_8753;
  assign x3159_0_io_sDone_1 = _T_8759;
  assign x3159_0_io_sDone_2 = _T_8765;
  assign x3159_0_io_w_0_addr_0 = x3297_wVec_0_addr_0;
  assign x3159_0_io_w_0_data = x3297_wVec_0_data;
  assign x3159_0_io_w_0_en = x3297_wVec_0_en;
  assign x3159_0_io_r_0_addr_0 = _T_8821_0_addr_0;
  assign x3159_0_io_r_0_en = _T_8821_0_en;
  assign x3159_0_io_r_1_addr_0 = _T_8821_1_addr_0;
  assign x3159_0_io_r_1_en = _T_8821_1_en;
  assign x3159_0_io_r_2_addr_0 = _T_8821_2_addr_0;
  assign x3159_0_io_r_2_en = _T_8821_2_en;
  assign x3159_0_io_r_3_addr_0 = _T_8821_3_addr_0;
  assign x3159_0_io_r_3_en = _T_8821_3_en;
  assign x3159_0_clock = clock;
  assign x3159_0_reset = reset;
  assign x3160_0_io_sEn_0 = x3428_base_en;
  assign x3160_0_io_sEn_1 = x3503_base_en;
  assign x3160_0_io_sDone_0 = _T_8771;
  assign x3160_0_io_sDone_1 = _T_8777;
  assign x3160_0_io_w_0_addr_0 = x3361_wVec_0_addr_0;
  assign x3160_0_io_w_0_data = x3361_wVec_0_data;
  assign x3160_0_io_w_0_en = x3361_wVec_0_en;
  assign x3160_0_io_r_0_addr_0 = _T_10136_0_addr_0;
  assign x3160_0_io_r_0_en = _T_10136_0_en;
  assign x3160_0_io_r_1_addr_0 = _T_10136_1_addr_0;
  assign x3160_0_io_r_1_en = _T_10136_1_en;
  assign x3160_0_io_r_2_addr_0 = _T_10136_2_addr_0;
  assign x3160_0_io_r_2_en = _T_10136_2_en;
  assign x3160_0_io_r_3_addr_0 = _T_10136_3_addr_0;
  assign x3160_0_io_r_3_en = _T_10136_3_en;
  assign x3160_0_clock = clock;
  assign x3160_0_reset = reset;
  assign x3161_0_io_sEn_0 = x3428_base_en;
  assign x3161_0_io_sEn_1 = x3503_base_en;
  assign x3161_0_io_sDone_0 = _T_8783;
  assign x3161_0_io_sDone_1 = _T_8789;
  assign x3161_0_io_w_0_addr_0 = x3424_wVec_0_addr_0;
  assign x3161_0_io_w_0_data = x3424_wVec_0_data;
  assign x3161_0_io_w_0_en = x3424_wVec_0_en;
  assign x3161_0_io_r_0_addr_0 = _T_8871_0_addr_0;
  assign x3161_0_io_r_0_en = _T_8871_0_en;
  assign x3161_0_io_r_1_addr_0 = _T_8871_1_addr_0;
  assign x3161_0_io_r_1_en = _T_8871_1_en;
  assign x3161_0_io_r_2_addr_0 = _T_8871_2_addr_0;
  assign x3161_0_io_r_2_en = _T_8871_2_en;
  assign x3161_0_io_r_3_addr_0 = _T_8871_3_addr_0;
  assign x3161_0_io_r_3_en = _T_8871_3_en;
  assign x3161_0_clock = clock;
  assign x3161_0_reset = reset;
  assign x3174_sm_io_input_enable = _T_2517;
  assign x3174_sm_io_input_stageDone_0 = x3167_done;
  assign x3174_sm_io_input_stageDone_1 = x3173_done;
  assign x3174_sm_io_input_stageMask_0 = x3167_mask;
  assign x3174_sm_io_input_stageMask_1 = x3173_mask;
  assign x3174_sm_io_input_rst = x3174_resetter;
  assign x3174_sm_clock = clock;
  assign x3174_sm_reset = reset;
  assign x3167_sm_io_input_enable = _T_8317;
  assign x3167_sm_io_input_ctr_done = _T_8351;
  assign x3167_sm_io_input_rst = x3167_resetter;
  assign x3167_sm_clock = clock;
  assign x3167_sm_reset = reset;
  assign x3173_sm_io_input_enable = _T_8363;
  assign x3173_sm_io_input_ctr_done = _T_8397;
  assign x3173_sm_io_input_rst = x3173_resetter;
  assign x3173_sm_clock = clock;
  assign x3173_sm_reset = reset;
  assign x3301_sm_io_input_enable = _T_2587;
  assign x3301_sm_io_input_stageDone_0 = x3237_done;
  assign x3301_sm_io_input_stageDone_1 = x3300_done;
  assign x3301_sm_io_input_stageMask_0 = x3237_mask;
  assign x3301_sm_io_input_stageMask_1 = x3300_mask;
  assign x3301_sm_io_input_rst = x3301_resetter;
  assign x3301_sm_clock = clock;
  assign x3301_sm_reset = reset;
  assign x3237_sm_io_input_enable = _T_2846;
  assign x3237_sm_io_input_stageDone_0 = x3208_done;
  assign x3237_sm_io_input_stageDone_1 = x3236_done;
  assign x3237_sm_io_input_stageMask_0 = x3208_mask;
  assign x3237_sm_io_input_stageMask_1 = x3236_mask;
  assign x3237_sm_io_input_rst = x3237_resetter;
  assign x3237_sm_clock = clock;
  assign x3237_sm_reset = reset;
  assign x3175_valid_srff_io_input_set = x3175_valid_options_0;
  assign x3175_valid_srff_io_input_reset = x3175_valid_stops_0;
  assign x3175_valid_srff_io_input_asyn_reset = _T_1601;
  assign x3175_valid_srff_clock = clock;
  assign x3175_valid_srff_reset = reset;
  assign x3176_io_in_0_data = _T_4485_0;
  assign x3176_io_in_0_en = _T_4499_0;
  assign x3176_io_deq_0 = _T_12077_0;
  assign x3176_clock = clock;
  assign x3176_reset = reset;
  assign x3208_sm_io_input_enable = _T_2984;
  assign x3208_sm_io_input_ctr_done = _T_3009;
  assign x3208_sm_io_input_rst = x3208_resetter;
  assign x3208_sm_clock = clock;
  assign x3208_sm_reset = reset;
  assign x3236_sm_io_input_enable = _T_3035;
  assign x3236_sm_io_input_stageDone_0 = x3220_done;
  assign x3236_sm_io_input_stageDone_1 = x3235_done;
  assign x3236_sm_io_input_stageMask_0 = x3220_mask;
  assign x3236_sm_io_input_stageMask_1 = x3235_mask;
  assign x3236_sm_io_input_rst = x3236_resetter;
  assign x3236_sm_clock = clock;
  assign x3236_sm_reset = reset;
  assign x3210_0_io_input_0_data = x3214_number;
  assign x3210_0_io_input_0_init = 32'h0;
  assign x3210_0_io_input_0_enable = _T_12093;
  assign x3210_0_io_input_0_reset = _T_12099;
  assign x3210_0_clock = clock;
  assign x3210_0_reset = reset;
  assign x3211_0_io_input_0_data = x3216_number;
  assign x3211_0_io_input_0_init = 32'h0;
  assign x3211_0_io_input_0_enable = _T_12093;
  assign x3211_0_io_input_0_reset = _T_12111;
  assign x3211_0_clock = clock;
  assign x3211_0_reset = reset;
  assign x3212_0_io_input_0_data = x3218_number;
  assign x3212_0_io_input_0_init = 32'h0;
  assign x3212_0_io_input_0_enable = _T_12093;
  assign x3212_0_io_input_0_reset = _T_12123;
  assign x3212_0_clock = clock;
  assign x3212_0_reset = reset;
  assign x3220_sm_io_input_enable = _T_3104;
  assign x3220_sm_io_input_ctr_done = _T_3127;
  assign x3220_sm_io_input_rst = x3220_resetter;
  assign x3220_sm_clock = clock;
  assign x3220_sm_reset = reset;
  assign x3223_io_input_stops_0 = _T_3139;
  assign x3223_io_input_reset = x3223_resetter;
  assign x3223_io_input_enable = x3223_en;
  assign x3223_clock = clock;
  assign x3223_reset = reset;
  assign x3235_sm_io_input_ctr_done = _T_3427;
  assign b1271 = _T_3531;
  assign x3300_sm_io_input_enable = _T_2915;
  assign x3300_sm_io_input_stageDone_0 = x3271_done;
  assign x3300_sm_io_input_stageDone_1 = x3299_done;
  assign x3300_sm_io_input_stageMask_0 = x3271_mask;
  assign x3300_sm_io_input_stageMask_1 = x3299_mask;
  assign x3300_sm_io_input_rst = x3300_resetter;
  assign x3300_sm_clock = clock;
  assign x3300_sm_reset = reset;
  assign x3238_valid_srff_io_input_set = x3238_valid_options_0;
  assign x3238_valid_srff_io_input_reset = x3238_valid_stops_0;
  assign x3238_valid_srff_io_input_asyn_reset = _T_1610;
  assign x3238_valid_srff_clock = clock;
  assign x3238_valid_srff_reset = reset;
  assign x3239_io_in_0_data = _T_7650_0;
  assign x3239_io_in_0_en = _T_7664_0;
  assign x3239_io_deq_0 = _T_11243_0;
  assign x3239_clock = clock;
  assign x3239_reset = reset;
  assign x3271_sm_io_input_enable = _T_4503;
  assign x3271_sm_io_input_ctr_done = _T_4528;
  assign x3271_sm_io_input_rst = x3271_resetter;
  assign x3271_sm_clock = clock;
  assign x3271_sm_reset = reset;
  assign x3299_sm_io_input_enable = _T_4554;
  assign x3299_sm_io_input_stageDone_0 = x3283_done;
  assign x3299_sm_io_input_stageDone_1 = x3298_done;
  assign x3299_sm_io_input_stageMask_0 = x3283_mask;
  assign x3299_sm_io_input_stageMask_1 = x3298_mask;
  assign x3299_sm_io_input_rst = x3299_resetter;
  assign x3299_sm_clock = clock;
  assign x3299_sm_reset = reset;
  assign x3273_0_io_input_0_data = x3277_number;
  assign x3273_0_io_input_0_init = 32'h0;
  assign x3273_0_io_input_0_enable = _T_11259;
  assign x3273_0_io_input_0_reset = _T_11265;
  assign x3273_0_clock = clock;
  assign x3273_0_reset = reset;
  assign x3274_0_io_input_0_data = x3279_number;
  assign x3274_0_io_input_0_init = 32'h0;
  assign x3274_0_io_input_0_enable = _T_11259;
  assign x3274_0_io_input_0_reset = _T_11277;
  assign x3274_0_clock = clock;
  assign x3274_0_reset = reset;
  assign x3275_0_io_input_0_data = x3281_number;
  assign x3275_0_io_input_0_init = 32'h0;
  assign x3275_0_io_input_0_enable = _T_11259;
  assign x3275_0_io_input_0_reset = _T_11289;
  assign x3275_0_clock = clock;
  assign x3275_0_reset = reset;
  assign x3283_sm_io_input_enable = _T_4623;
  assign x3283_sm_io_input_ctr_done = _T_4646;
  assign x3283_sm_io_input_rst = x3283_resetter;
  assign x3283_sm_clock = clock;
  assign x3283_sm_reset = reset;
  assign x3286_io_input_stops_0 = _T_4658;
  assign x3286_io_input_reset = x3286_resetter;
  assign x3286_io_input_enable = x3286_en;
  assign x3286_clock = clock;
  assign x3286_reset = reset;
  assign x3298_sm_io_input_ctr_done = _T_4946;
  assign b1332 = _T_5050;
  assign x3428_sm_io_input_enable = _T_2657;
  assign x3428_sm_io_input_stageDone_0 = x3364_done;
  assign x3428_sm_io_input_stageDone_1 = x3427_done;
  assign x3428_sm_io_input_stageMask_0 = x3364_mask;
  assign x3428_sm_io_input_stageMask_1 = x3427_mask;
  assign x3428_sm_io_input_rst = x3428_resetter;
  assign x3428_sm_clock = clock;
  assign x3428_sm_reset = reset;
  assign x3364_sm_io_input_enable = _T_3596;
  assign x3364_sm_io_input_stageDone_0 = x3335_done;
  assign x3364_sm_io_input_stageDone_1 = x3363_done;
  assign x3364_sm_io_input_stageMask_0 = x3335_mask;
  assign x3364_sm_io_input_stageMask_1 = x3363_mask;
  assign x3364_sm_io_input_rst = x3364_resetter;
  assign x3364_sm_clock = clock;
  assign x3364_sm_reset = reset;
  assign x3302_valid_srff_io_input_set = x3302_valid_options_0;
  assign x3302_valid_srff_io_input_reset = x3302_valid_stops_0;
  assign x3302_valid_srff_io_input_asyn_reset = _T_1619;
  assign x3302_valid_srff_clock = clock;
  assign x3302_valid_srff_reset = reset;
  assign x3303_io_in_0_data = _T_11214_0;
  assign x3303_io_in_0_en = _T_11228_0;
  assign x3303_io_deq_0 = _T_12385_0;
  assign x3303_clock = clock;
  assign x3303_reset = reset;
  assign x3335_sm_io_input_enable = _T_9318;
  assign x3335_sm_io_input_ctr_done = _T_9343;
  assign x3335_sm_io_input_rst = x3335_resetter;
  assign x3335_sm_clock = clock;
  assign x3335_sm_reset = reset;
  assign x3363_sm_io_input_enable = _T_9369;
  assign x3363_sm_io_input_stageDone_0 = x3347_done;
  assign x3363_sm_io_input_stageDone_1 = x3362_done;
  assign x3363_sm_io_input_stageMask_0 = x3347_mask;
  assign x3363_sm_io_input_stageMask_1 = x3362_mask;
  assign x3363_sm_io_input_rst = x3363_resetter;
  assign x3363_sm_clock = clock;
  assign x3363_sm_reset = reset;
  assign x3337_0_io_input_0_data = x3341_number;
  assign x3337_0_io_input_0_init = 32'h0;
  assign x3337_0_io_input_0_enable = _T_12401;
  assign x3337_0_io_input_0_reset = _T_12407;
  assign x3337_0_clock = clock;
  assign x3337_0_reset = reset;
  assign x3338_0_io_input_0_data = x3343_number;
  assign x3338_0_io_input_0_init = 32'h0;
  assign x3338_0_io_input_0_enable = _T_12401;
  assign x3338_0_io_input_0_reset = _T_12419;
  assign x3338_0_clock = clock;
  assign x3338_0_reset = reset;
  assign x3339_0_io_input_0_data = x3345_number;
  assign x3339_0_io_input_0_init = 32'h0;
  assign x3339_0_io_input_0_enable = _T_12401;
  assign x3339_0_io_input_0_reset = _T_12431;
  assign x3339_0_clock = clock;
  assign x3339_0_reset = reset;
  assign x3347_sm_io_input_enable = _T_9438;
  assign x3347_sm_io_input_ctr_done = _T_9461;
  assign x3347_sm_io_input_rst = x3347_resetter;
  assign x3347_sm_clock = clock;
  assign x3347_sm_reset = reset;
  assign x3350_io_input_stops_0 = _T_9473;
  assign x3350_io_input_reset = x3350_resetter;
  assign x3350_io_input_enable = x3350_en;
  assign x3350_clock = clock;
  assign x3350_reset = reset;
  assign x3362_sm_io_input_ctr_done = _T_9761;
  assign b1394 = _T_9865;
  assign x3427_sm_io_input_enable = _T_3665;
  assign x3427_sm_io_input_stageDone_0 = x3398_done;
  assign x3427_sm_io_input_stageDone_1 = x3426_done;
  assign x3427_sm_io_input_stageMask_0 = x3398_mask;
  assign x3427_sm_io_input_stageMask_1 = x3426_mask;
  assign x3427_sm_io_input_rst = x3427_resetter;
  assign x3427_sm_clock = clock;
  assign x3427_sm_reset = reset;
  assign x3365_valid_srff_io_input_set = x3365_valid_options_0;
  assign x3365_valid_srff_io_input_reset = x3365_valid_stops_0;
  assign x3365_valid_srff_io_input_asyn_reset = _T_1628;
  assign x3365_valid_srff_clock = clock;
  assign x3365_valid_srff_reset = reset;
  assign x3366_io_in_0_data = _T_8299_0;
  assign x3366_io_in_0_en = _T_8313_0;
  assign x3366_io_deq_0 = _T_12443_0;
  assign x3366_clock = clock;
  assign x3366_reset = reset;
  assign x3398_sm_io_input_enable = _T_3734;
  assign x3398_sm_io_input_ctr_done = _T_3759;
  assign x3398_sm_io_input_rst = x3398_resetter;
  assign x3398_sm_clock = clock;
  assign x3398_sm_reset = reset;
  assign x3426_sm_io_input_enable = _T_3785;
  assign x3426_sm_io_input_stageDone_0 = x3410_done;
  assign x3426_sm_io_input_stageDone_1 = x3425_done;
  assign x3426_sm_io_input_stageMask_0 = x3410_mask;
  assign x3426_sm_io_input_stageMask_1 = x3425_mask;
  assign x3426_sm_io_input_rst = x3426_resetter;
  assign x3426_sm_clock = clock;
  assign x3426_sm_reset = reset;
  assign x3400_0_io_input_0_data = x3404_number;
  assign x3400_0_io_input_0_init = 32'h0;
  assign x3400_0_io_input_0_enable = _T_12459;
  assign x3400_0_io_input_0_reset = _T_12465;
  assign x3400_0_clock = clock;
  assign x3400_0_reset = reset;
  assign x3401_0_io_input_0_data = x3406_number;
  assign x3401_0_io_input_0_init = 32'h0;
  assign x3401_0_io_input_0_enable = _T_12459;
  assign x3401_0_io_input_0_reset = _T_12477;
  assign x3401_0_clock = clock;
  assign x3401_0_reset = reset;
  assign x3402_0_io_input_0_data = x3408_number;
  assign x3402_0_io_input_0_init = 32'h0;
  assign x3402_0_io_input_0_enable = _T_12459;
  assign x3402_0_io_input_0_reset = _T_12489;
  assign x3402_0_clock = clock;
  assign x3402_0_reset = reset;
  assign x3410_sm_io_input_enable = _T_11449;
  assign x3410_sm_io_input_ctr_done = _T_11472;
  assign x3410_sm_io_input_rst = x3410_resetter;
  assign x3410_sm_clock = clock;
  assign x3410_sm_reset = reset;
  assign x3413_io_input_stops_0 = _T_11484;
  assign x3413_io_input_reset = x3413_resetter;
  assign x3413_io_input_enable = x3413_en;
  assign x3413_clock = clock;
  assign x3413_reset = reset;
  assign x3425_sm_io_input_ctr_done = _T_11772;
  assign b1455 = _T_11876;
  assign x3429_0_io_input_next = x3464_number;
  assign x3429_0_io_input_enable = _T_10565;
  assign x3429_0_io_input_reset = _T_10569;
  assign x3429_0_clock = clock;
  assign x3429_0_reset = reset;
  assign x3429_1_io_sEn_0 = x3503_base_en;
  assign x3429_1_io_sEn_1 = x3514_base_en;
  assign x3429_1_io_sDone_0 = _T_8711;
  assign x3429_1_io_sDone_1 = _T_8717;
  assign x3429_1_io_input_0_data = x3465_number;
  assign x3429_1_io_input_0_enable = _T_10577;
  assign x3429_1_io_input_0_reset = _T_10581;
  assign x3429_1_clock = clock;
  assign x3429_1_reset = reset;
  assign x3430_0_io_input_next = x3500_number;
  assign x3430_0_io_input_enable = _T_9300;
  assign x3430_0_io_input_reset = _T_9304;
  assign x3430_0_clock = clock;
  assign x3430_0_reset = reset;
  assign x3430_1_io_sEn_0 = x3503_base_en;
  assign x3430_1_io_sEn_1 = x3514_base_en;
  assign x3430_1_io_sDone_0 = _T_8723;
  assign x3430_1_io_sDone_1 = _T_8729;
  assign x3430_1_io_input_0_data = x3501_number;
  assign x3430_1_io_input_0_enable = _T_9312;
  assign x3430_1_io_input_0_reset = _T_9316;
  assign x3430_1_clock = clock;
  assign x3430_1_reset = reset;
  assign x3503_sm_io_input_enable = _T_2729;
  assign x3503_sm_io_input_stageDone_0 = x3466_done;
  assign x3503_sm_io_input_stageDone_1 = x3502_done;
  assign x3503_sm_io_input_stageMask_0 = x3466_mask;
  assign x3503_sm_io_input_stageMask_1 = x3502_mask;
  assign x3503_sm_io_input_rst = x3503_resetter;
  assign x3503_sm_clock = clock;
  assign x3503_sm_reset = reset;
  assign x3433_io_input_stops_0 = _T_5115;
  assign x3433_io_input_reset = x3433_resetter;
  assign x3433_io_input_enable = x3433_en;
  assign x3433_clock = clock;
  assign x3433_reset = reset;
  assign x3466_sm_io_input_enable = _T_5382;
  assign x3466_sm_io_input_ctr_done = _T_5409;
  assign x3466_sm_io_input_rst = x3466_resetter;
  assign x3466_sm_clock = clock;
  assign x3466_sm_reset = reset;
  assign b1483 = _T_5518;
  assign b1484 = _T_5648;
  assign b1485 = _T_5778;
  assign b1486 = _T_5908;
  assign x3469_io_input_stops_0 = _T_5973;
  assign x3469_io_input_reset = x3469_resetter;
  assign x3469_io_input_enable = x3469_en;
  assign x3469_clock = clock;
  assign x3469_reset = reset;
  assign x3502_sm_io_input_enable = _T_6240;
  assign x3502_sm_io_input_ctr_done = _T_6267;
  assign x3502_sm_io_input_rst = x3502_resetter;
  assign x3502_sm_clock = clock;
  assign x3502_sm_reset = reset;
  assign b1524 = _T_6376;
  assign b1525 = _T_6506;
  assign b1526 = _T_6636;
  assign b1527 = _T_6766;
  assign x3514_sm_io_input_enable = _T_2799;
  assign x3514_sm_io_input_ctr_done = _T_2833;
  assign x3514_sm_io_input_rst = x3514_resetter;
  assign x3514_sm_clock = clock;
  assign x3514_sm_reset = reset;
  assign b1204_chain_io_sEn_0 = x3174_en;
  assign b1204_chain_io_sEn_1 = x3301_en;
  assign b1204_chain_io_sEn_2 = x3428_en;
  assign b1204_chain_io_sEn_3 = x3503_en;
  assign b1204_chain_io_sEn_4 = x3514_en;
  assign b1204_chain_io_sDone_0 = _T_8573;
  assign b1204_chain_io_sDone_1 = _T_8579;
  assign b1204_chain_io_sDone_2 = _T_8585;
  assign b1204_chain_io_sDone_3 = _T_8591;
  assign b1204_chain_io_sDone_4 = _T_8597;
  assign b1204_chain_io_input_0_data = b1204;
  assign b1204_chain_io_input_0_enable = x3515_sm_io_output_ctr_inc;
  assign b1204_chain_io_input_0_reset = _T_2136;
  assign b1204_chain_clock = clock;
  assign b1204_chain_reset = reset;
  assign b1205_chain_io_sEn_0 = x3174_en;
  assign b1205_chain_io_sEn_1 = x3301_en;
  assign b1205_chain_io_sEn_2 = x3428_en;
  assign b1205_chain_io_sEn_3 = x3503_en;
  assign b1205_chain_io_sEn_4 = x3514_en;
  assign b1205_chain_io_sDone_0 = _T_8603;
  assign b1205_chain_io_sDone_1 = _T_8609;
  assign b1205_chain_io_sDone_2 = _T_8615;
  assign b1205_chain_io_sDone_3 = _T_8621;
  assign b1205_chain_io_sDone_4 = _T_8627;
  assign b1205_chain_io_input_0_data = b1205;
  assign b1205_chain_io_input_0_enable = x3515_sm_io_output_ctr_inc;
  assign b1205_chain_io_input_0_reset = _T_2273;
  assign b1205_chain_clock = clock;
  assign b1205_chain_reset = reset;
  assign x3518_sm_io_input_enable = _T_2426;
  assign x3518_sm_io_input_ctr_done = _T_2460;
  assign x3518_sm_io_input_rst = x3518_resetter;
  assign x3518_sm_clock = clock;
  assign x3518_sm_reset = reset;
  assign RetimeWrapper_1_io_flow = 1'h1;
  assign RetimeWrapper_1_io_in = reset;
  assign RetimeWrapper_1_clock = clock;
  assign RetimeWrapper_1_reset = reset;
  assign _T_1702 = RetimeWrapper_1_io_out;
  assign retime_counter_io_input_reset = reset;
  assign retime_counter_clock = clock;
  assign retime_counter_reset = reset;
  assign RetimeWrapper_2_io_flow = 1'h1;
  assign RetimeWrapper_2_io_in = retime_counter_io_output_done;
  assign RetimeWrapper_2_clock = clock;
  assign RetimeWrapper_2_reset = reset;
  assign _T_1710 = RetimeWrapper_2_io_out;
  assign _T_1722_number = _T_1755;
  assign _T_1724_number = _T_1734;
  assign _T_1734 = _T_1739;
  assign x35150_range_number = _T_1770;
  assign _T_1770 = _T_1774;
  assign x35150_hops_number = _T_1786_number;
  assign _T_1786_number = _T_1796;
  assign _T_1788_number = _T_1784[31:0];
  assign _T_1796 = _T_1788_number;
  assign _T_1805_number = {{32'd0}, _T_1806};
  assign x35150_leftover_number = _T_1815;
  assign _T_1815 = _T_1881;
  assign _T_1909_number = _T_1919;
  assign _T_1911_number = x35150_adjustment;
  assign _T_1919 = _T_1928;
  assign _T_1930_number = _T_1962;
  assign _T_1932_number = _T_1942;
  assign _T_1934_number = _T_1955;
  assign _T_1942 = _T_1947;
  assign _T_1955 = _T_1960;
  assign _T_1964_number = _T_1972;
  assign _T_1972 = _T_1976;
  assign _T_2075_number = _T_2085;
  assign _T_2077_number = _T_2096;
  assign _T_2085 = b1202_number;
  assign _T_2096 = x3153_number;
  assign RetimeWrapper_3_io_flow = 1'h1;
  assign RetimeWrapper_3_io_in = b1204_chain_reset;
  assign RetimeWrapper_3_clock = clock;
  assign RetimeWrapper_3_reset = reset;
  assign _T_2136 = RetimeWrapper_3_io_out;
  assign _T_2212_number = _T_2222;
  assign _T_2214_number = _T_2233;
  assign _T_2222 = b1203_number;
  assign _T_2233 = x3153_number;
  assign RetimeWrapper_4_io_flow = 1'h1;
  assign RetimeWrapper_4_io_in = b1205_chain_reset;
  assign RetimeWrapper_4_clock = clock;
  assign RetimeWrapper_4_reset = reset;
  assign _T_2273 = RetimeWrapper_4_io_out;
  assign RetimeWrapper_5_io_flow = 1'h1;
  assign RetimeWrapper_5_io_in = x3515_sm_io_output_stageEnable_0;
  assign RetimeWrapper_5_clock = clock;
  assign RetimeWrapper_5_reset = reset;
  assign _T_2280 = RetimeWrapper_5_io_out;
  assign RetimeWrapper_6_io_flow = 1'h1;
  assign RetimeWrapper_6_io_in = _T_2283;
  assign RetimeWrapper_6_clock = clock;
  assign RetimeWrapper_6_reset = reset;
  assign _T_2287 = RetimeWrapper_6_io_out;
  assign RetimeWrapper_7_io_flow = 1'h1;
  assign RetimeWrapper_7_io_in = x3515_sm_io_output_rst_en;
  assign RetimeWrapper_7_clock = clock;
  assign RetimeWrapper_7_reset = reset;
  assign _T_2294 = RetimeWrapper_7_io_out;
  assign RetimeWrapper_8_io_flow = 1'h1;
  assign RetimeWrapper_8_io_in = x3515_sm_io_output_stageEnable_1;
  assign RetimeWrapper_8_clock = clock;
  assign RetimeWrapper_8_reset = reset;
  assign _T_2300 = RetimeWrapper_8_io_out;
  assign RetimeWrapper_9_io_flow = 1'h1;
  assign RetimeWrapper_9_io_in = _T_2303;
  assign RetimeWrapper_9_clock = clock;
  assign RetimeWrapper_9_reset = reset;
  assign _T_2307 = RetimeWrapper_9_io_out;
  assign RetimeWrapper_10_io_flow = 1'h1;
  assign RetimeWrapper_10_io_in = x3515_sm_io_output_rst_en;
  assign RetimeWrapper_10_clock = clock;
  assign RetimeWrapper_10_reset = reset;
  assign _T_2314 = RetimeWrapper_10_io_out;
  assign RetimeWrapper_11_io_flow = 1'h1;
  assign RetimeWrapper_11_io_in = x3515_sm_io_output_stageEnable_2;
  assign RetimeWrapper_11_clock = clock;
  assign RetimeWrapper_11_reset = reset;
  assign _T_2320 = RetimeWrapper_11_io_out;
  assign RetimeWrapper_12_io_flow = 1'h1;
  assign RetimeWrapper_12_io_in = _T_2323;
  assign RetimeWrapper_12_clock = clock;
  assign RetimeWrapper_12_reset = reset;
  assign _T_2327 = RetimeWrapper_12_io_out;
  assign RetimeWrapper_13_io_flow = 1'h1;
  assign RetimeWrapper_13_io_in = x3515_sm_io_output_rst_en;
  assign RetimeWrapper_13_clock = clock;
  assign RetimeWrapper_13_reset = reset;
  assign _T_2334 = RetimeWrapper_13_io_out;
  assign RetimeWrapper_14_io_flow = 1'h1;
  assign RetimeWrapper_14_io_in = x3515_sm_io_output_stageEnable_3;
  assign RetimeWrapper_14_clock = clock;
  assign RetimeWrapper_14_reset = reset;
  assign _T_2340 = RetimeWrapper_14_io_out;
  assign RetimeWrapper_15_io_flow = 1'h1;
  assign RetimeWrapper_15_io_in = _T_2343;
  assign RetimeWrapper_15_clock = clock;
  assign RetimeWrapper_15_reset = reset;
  assign _T_2347 = RetimeWrapper_15_io_out;
  assign RetimeWrapper_16_io_flow = 1'h1;
  assign RetimeWrapper_16_io_in = x3515_sm_io_output_rst_en;
  assign RetimeWrapper_16_clock = clock;
  assign RetimeWrapper_16_reset = reset;
  assign _T_2354 = RetimeWrapper_16_io_out;
  assign RetimeWrapper_17_io_flow = 1'h1;
  assign RetimeWrapper_17_io_in = x3515_sm_io_output_stageEnable_4;
  assign RetimeWrapper_17_clock = clock;
  assign RetimeWrapper_17_reset = reset;
  assign _T_2360 = RetimeWrapper_17_io_out;
  assign RetimeWrapper_18_io_flow = 1'h1;
  assign RetimeWrapper_18_io_in = _T_2363;
  assign RetimeWrapper_18_clock = clock;
  assign RetimeWrapper_18_reset = reset;
  assign _T_2367 = RetimeWrapper_18_io_out;
  assign RetimeWrapper_19_io_flow = 1'h1;
  assign RetimeWrapper_19_io_in = x3515_sm_io_output_rst_en;
  assign RetimeWrapper_19_clock = clock;
  assign RetimeWrapper_19_reset = reset;
  assign _T_2374 = RetimeWrapper_19_io_out;
  assign RetimeWrapper_20_io_flow = 1'h1;
  assign RetimeWrapper_20_io_in = b1202_chain_reset;
  assign RetimeWrapper_20_clock = clock;
  assign RetimeWrapper_20_reset = reset;
  assign _T_2380 = RetimeWrapper_20_io_out;
  assign RetimeWrapper_21_io_flow = 1'h1;
  assign RetimeWrapper_21_io_in = b1203_chain_reset;
  assign RetimeWrapper_21_clock = clock;
  assign RetimeWrapper_21_reset = reset;
  assign _T_2387 = RetimeWrapper_21_io_out;
  assign RetimeWrapper_22_io_flow = 1'h1;
  assign RetimeWrapper_22_io_in = 1'h0;
  assign RetimeWrapper_22_clock = clock;
  assign RetimeWrapper_22_reset = reset;
  assign _T_2394 = RetimeWrapper_22_io_out;
  assign _T_2398_number = _T_2408;
  assign _T_2408 = x3153_number;
  assign RetimeWrapper_23_io_flow = 1'h1;
  assign RetimeWrapper_23_io_in = _T_2454;
  assign RetimeWrapper_23_clock = clock;
  assign RetimeWrapper_23_reset = reset;
  assign _T_2458 = RetimeWrapper_23_io_out;
  assign RetimeWrapper_24_io_flow = 1'h1;
  assign RetimeWrapper_24_io_in = 1'h0;
  assign RetimeWrapper_24_clock = clock;
  assign RetimeWrapper_24_reset = reset;
  assign _T_2466 = RetimeWrapper_24_io_out;
  assign RetimeWrapper_25_io_flow = 1'h1;
  assign RetimeWrapper_25_io_in = RootController_sm_io_output_stageEnable_0;
  assign RetimeWrapper_25_clock = clock;
  assign RetimeWrapper_25_reset = reset;
  assign _T_2476 = RetimeWrapper_25_io_out;
  assign RetimeWrapper_26_io_flow = 1'h1;
  assign RetimeWrapper_26_io_in = _T_1992;
  assign RetimeWrapper_26_clock = clock;
  assign RetimeWrapper_26_reset = reset;
  assign _T_2483 = RetimeWrapper_26_io_out;
  assign RetimeWrapper_27_io_flow = 1'h1;
  assign RetimeWrapper_27_io_in = RootController_sm_io_output_rst_en;
  assign RetimeWrapper_27_clock = clock;
  assign RetimeWrapper_27_reset = reset;
  assign _T_2490 = RetimeWrapper_27_io_out;
  assign RetimeWrapper_28_io_flow = 1'h1;
  assign RetimeWrapper_28_io_in = RootController_sm_io_output_stageEnable_1;
  assign RetimeWrapper_28_clock = clock;
  assign RetimeWrapper_28_reset = reset;
  assign _T_2496 = RetimeWrapper_28_io_out;
  assign RetimeWrapper_29_io_flow = 1'h1;
  assign RetimeWrapper_29_io_in = _T_2441;
  assign RetimeWrapper_29_clock = clock;
  assign RetimeWrapper_29_reset = reset;
  assign _T_2503 = RetimeWrapper_29_io_out;
  assign RetimeWrapper_30_io_flow = 1'h1;
  assign RetimeWrapper_30_io_in = RootController_sm_io_output_rst_en;
  assign RetimeWrapper_30_clock = clock;
  assign RetimeWrapper_30_reset = reset;
  assign _T_2510 = RetimeWrapper_30_io_out;
  assign done_latch_io_input_set = RootController_done;
  assign done_latch_io_input_reset = RootController_resetter;
  assign done_latch_io_input_asyn_reset = RootController_resetter;
  assign done_latch_clock = clock;
  assign done_latch_reset = reset;
  assign RetimeWrapper_31_io_flow = 1'h1;
  assign RetimeWrapper_31_io_in = x3515_ctr_trivial;
  assign RetimeWrapper_31_clock = clock;
  assign RetimeWrapper_31_reset = reset;
  assign _T_2541 = RetimeWrapper_31_io_out;
  assign RetimeWrapper_32_io_flow = 1'h1;
  assign RetimeWrapper_32_io_in = x3174_sm_io_output_stageEnable_0;
  assign RetimeWrapper_32_clock = clock;
  assign RetimeWrapper_32_reset = reset;
  assign _T_2549 = RetimeWrapper_32_io_out;
  assign RetimeWrapper_33_io_flow = 1'h1;
  assign RetimeWrapper_33_io_in = _T_2552;
  assign RetimeWrapper_33_clock = clock;
  assign RetimeWrapper_33_reset = reset;
  assign _T_2556 = RetimeWrapper_33_io_out;
  assign RetimeWrapper_34_io_flow = 1'h1;
  assign RetimeWrapper_34_io_in = x3174_sm_io_output_rst_en;
  assign RetimeWrapper_34_clock = clock;
  assign RetimeWrapper_34_reset = reset;
  assign _T_2563 = RetimeWrapper_34_io_out;
  assign RetimeWrapper_35_io_flow = 1'h1;
  assign RetimeWrapper_35_io_in = x3174_sm_io_output_stageEnable_1;
  assign RetimeWrapper_35_clock = clock;
  assign RetimeWrapper_35_reset = reset;
  assign _T_2569 = RetimeWrapper_35_io_out;
  assign RetimeWrapper_36_io_flow = 1'h1;
  assign RetimeWrapper_36_io_in = _T_2572;
  assign RetimeWrapper_36_clock = clock;
  assign RetimeWrapper_36_reset = reset;
  assign _T_2576 = RetimeWrapper_36_io_out;
  assign RetimeWrapper_37_io_flow = 1'h1;
  assign RetimeWrapper_37_io_in = x3174_sm_io_output_rst_en;
  assign RetimeWrapper_37_clock = clock;
  assign RetimeWrapper_37_reset = reset;
  assign _T_2583 = RetimeWrapper_37_io_out;
  assign RetimeWrapper_38_io_flow = 1'h1;
  assign RetimeWrapper_38_io_in = x3515_ctr_trivial;
  assign RetimeWrapper_38_clock = clock;
  assign RetimeWrapper_38_reset = reset;
  assign _T_2611 = RetimeWrapper_38_io_out;
  assign RetimeWrapper_39_io_flow = 1'h1;
  assign RetimeWrapper_39_io_in = x3301_sm_io_output_stageEnable_0;
  assign RetimeWrapper_39_clock = clock;
  assign RetimeWrapper_39_reset = reset;
  assign _T_2619 = RetimeWrapper_39_io_out;
  assign RetimeWrapper_40_io_flow = 1'h1;
  assign RetimeWrapper_40_io_in = _T_2622;
  assign RetimeWrapper_40_clock = clock;
  assign RetimeWrapper_40_reset = reset;
  assign _T_2626 = RetimeWrapper_40_io_out;
  assign RetimeWrapper_41_io_flow = 1'h1;
  assign RetimeWrapper_41_io_in = x3301_sm_io_output_rst_en;
  assign RetimeWrapper_41_clock = clock;
  assign RetimeWrapper_41_reset = reset;
  assign _T_2633 = RetimeWrapper_41_io_out;
  assign RetimeWrapper_42_io_flow = 1'h1;
  assign RetimeWrapper_42_io_in = x3301_sm_io_output_stageEnable_1;
  assign RetimeWrapper_42_clock = clock;
  assign RetimeWrapper_42_reset = reset;
  assign _T_2639 = RetimeWrapper_42_io_out;
  assign RetimeWrapper_43_io_flow = 1'h1;
  assign RetimeWrapper_43_io_in = _T_2642;
  assign RetimeWrapper_43_clock = clock;
  assign RetimeWrapper_43_reset = reset;
  assign _T_2646 = RetimeWrapper_43_io_out;
  assign RetimeWrapper_44_io_flow = 1'h1;
  assign RetimeWrapper_44_io_in = x3301_sm_io_output_rst_en;
  assign RetimeWrapper_44_clock = clock;
  assign RetimeWrapper_44_reset = reset;
  assign _T_2653 = RetimeWrapper_44_io_out;
  assign RetimeWrapper_45_io_flow = 1'h1;
  assign RetimeWrapper_45_io_in = x3515_ctr_trivial;
  assign RetimeWrapper_45_clock = clock;
  assign RetimeWrapper_45_reset = reset;
  assign _T_2681 = RetimeWrapper_45_io_out;
  assign RetimeWrapper_46_io_flow = 1'h1;
  assign RetimeWrapper_46_io_in = x3428_sm_io_output_stageEnable_0;
  assign RetimeWrapper_46_clock = clock;
  assign RetimeWrapper_46_reset = reset;
  assign _T_2689 = RetimeWrapper_46_io_out;
  assign RetimeWrapper_47_io_flow = 1'h1;
  assign RetimeWrapper_47_io_in = _T_2692;
  assign RetimeWrapper_47_clock = clock;
  assign RetimeWrapper_47_reset = reset;
  assign _T_2696 = RetimeWrapper_47_io_out;
  assign RetimeWrapper_48_io_flow = 1'h1;
  assign RetimeWrapper_48_io_in = x3428_sm_io_output_rst_en;
  assign RetimeWrapper_48_clock = clock;
  assign RetimeWrapper_48_reset = reset;
  assign _T_2703 = RetimeWrapper_48_io_out;
  assign RetimeWrapper_49_io_flow = 1'h1;
  assign RetimeWrapper_49_io_in = x3428_sm_io_output_stageEnable_1;
  assign RetimeWrapper_49_clock = clock;
  assign RetimeWrapper_49_reset = reset;
  assign _T_2709 = RetimeWrapper_49_io_out;
  assign RetimeWrapper_50_io_flow = 1'h1;
  assign RetimeWrapper_50_io_in = _T_2712;
  assign RetimeWrapper_50_clock = clock;
  assign RetimeWrapper_50_reset = reset;
  assign _T_2716 = RetimeWrapper_50_io_out;
  assign RetimeWrapper_51_io_flow = 1'h1;
  assign RetimeWrapper_51_io_in = x3428_sm_io_output_rst_en;
  assign RetimeWrapper_51_clock = clock;
  assign RetimeWrapper_51_reset = reset;
  assign _T_2723 = RetimeWrapper_51_io_out;
  assign RetimeWrapper_52_io_flow = 1'h1;
  assign RetimeWrapper_52_io_in = x3515_ctr_trivial;
  assign RetimeWrapper_52_clock = clock;
  assign RetimeWrapper_52_reset = reset;
  assign _T_2753 = RetimeWrapper_52_io_out;
  assign RetimeWrapper_53_io_flow = 1'h1;
  assign RetimeWrapper_53_io_in = x3503_sm_io_output_stageEnable_0;
  assign RetimeWrapper_53_clock = clock;
  assign RetimeWrapper_53_reset = reset;
  assign _T_2761 = RetimeWrapper_53_io_out;
  assign RetimeWrapper_54_io_flow = 1'h1;
  assign RetimeWrapper_54_io_in = _T_2764;
  assign RetimeWrapper_54_clock = clock;
  assign RetimeWrapper_54_reset = reset;
  assign _T_2768 = RetimeWrapper_54_io_out;
  assign RetimeWrapper_55_io_flow = 1'h1;
  assign RetimeWrapper_55_io_in = x3503_sm_io_output_rst_en;
  assign RetimeWrapper_55_clock = clock;
  assign RetimeWrapper_55_reset = reset;
  assign _T_2775 = RetimeWrapper_55_io_out;
  assign RetimeWrapper_56_io_flow = 1'h1;
  assign RetimeWrapper_56_io_in = x3503_sm_io_output_stageEnable_1;
  assign RetimeWrapper_56_clock = clock;
  assign RetimeWrapper_56_reset = reset;
  assign _T_2781 = RetimeWrapper_56_io_out;
  assign RetimeWrapper_57_io_flow = 1'h1;
  assign RetimeWrapper_57_io_in = _T_2784;
  assign RetimeWrapper_57_clock = clock;
  assign RetimeWrapper_57_reset = reset;
  assign _T_2788 = RetimeWrapper_57_io_out;
  assign RetimeWrapper_58_io_flow = 1'h1;
  assign RetimeWrapper_58_io_in = x3503_sm_io_output_rst_en;
  assign RetimeWrapper_58_clock = clock;
  assign RetimeWrapper_58_reset = reset;
  assign _T_2795 = RetimeWrapper_58_io_out;
  assign RetimeWrapper_59_io_flow = 1'h1;
  assign RetimeWrapper_59_io_in = _T_2827;
  assign RetimeWrapper_59_clock = clock;
  assign RetimeWrapper_59_reset = reset;
  assign _T_2831 = RetimeWrapper_59_io_out;
  assign RetimeWrapper_60_io_flow = 1'h1;
  assign RetimeWrapper_60_io_in = x3515_ctr_trivial;
  assign RetimeWrapper_60_clock = clock;
  assign RetimeWrapper_60_reset = reset;
  assign RetimeWrapper_61_io_flow = 1'h1;
  assign RetimeWrapper_61_io_in = x3301_ctr_trivial;
  assign RetimeWrapper_61_clock = clock;
  assign RetimeWrapper_61_reset = reset;
  assign _T_2859 = RetimeWrapper_61_io_out;
  assign RetimeWrapper_62_io_flow = 1'h1;
  assign RetimeWrapper_62_io_in = x3237_sm_io_output_stageEnable_0;
  assign RetimeWrapper_62_clock = clock;
  assign RetimeWrapper_62_reset = reset;
  assign _T_2867 = RetimeWrapper_62_io_out;
  assign RetimeWrapper_63_io_flow = 1'h1;
  assign RetimeWrapper_63_io_in = _T_2870;
  assign RetimeWrapper_63_clock = clock;
  assign RetimeWrapper_63_reset = reset;
  assign _T_2874 = RetimeWrapper_63_io_out;
  assign RetimeWrapper_64_io_flow = 1'h1;
  assign RetimeWrapper_64_io_in = _T_2879;
  assign RetimeWrapper_64_clock = clock;
  assign RetimeWrapper_64_reset = reset;
  assign _T_2883 = RetimeWrapper_64_io_out;
  assign RetimeWrapper_65_io_flow = 1'h1;
  assign RetimeWrapper_65_io_in = x3237_sm_io_output_rst_en;
  assign RetimeWrapper_65_clock = clock;
  assign RetimeWrapper_65_reset = reset;
  assign _T_2892 = RetimeWrapper_65_io_out;
  assign RetimeWrapper_66_io_flow = 1'h1;
  assign RetimeWrapper_66_io_in = x3237_sm_io_output_stageEnable_1;
  assign RetimeWrapper_66_clock = clock;
  assign RetimeWrapper_66_reset = reset;
  assign _T_2898 = RetimeWrapper_66_io_out;
  assign RetimeWrapper_67_io_flow = 1'h1;
  assign RetimeWrapper_67_io_in = _T_2901;
  assign RetimeWrapper_67_clock = clock;
  assign RetimeWrapper_67_reset = reset;
  assign _T_2905 = RetimeWrapper_67_io_out;
  assign RetimeWrapper_68_io_flow = 1'h1;
  assign RetimeWrapper_68_io_in = x3237_sm_io_output_rst_en;
  assign RetimeWrapper_68_clock = clock;
  assign RetimeWrapper_68_reset = reset;
  assign _T_2912 = RetimeWrapper_68_io_out;
  assign RetimeWrapper_69_io_flow = 1'h1;
  assign RetimeWrapper_69_io_in = x3301_ctr_trivial;
  assign RetimeWrapper_69_clock = clock;
  assign RetimeWrapper_69_reset = reset;
  assign _T_2928 = RetimeWrapper_69_io_out;
  assign RetimeWrapper_70_io_flow = 1'h1;
  assign RetimeWrapper_70_io_in = x3300_sm_io_output_stageEnable_0;
  assign RetimeWrapper_70_clock = clock;
  assign RetimeWrapper_70_reset = reset;
  assign _T_2936 = RetimeWrapper_70_io_out;
  assign RetimeWrapper_71_io_flow = 1'h1;
  assign RetimeWrapper_71_io_in = _T_2939;
  assign RetimeWrapper_71_clock = clock;
  assign RetimeWrapper_71_reset = reset;
  assign _T_2943 = RetimeWrapper_71_io_out;
  assign RetimeWrapper_72_io_flow = 1'h1;
  assign RetimeWrapper_72_io_in = _T_2948;
  assign RetimeWrapper_72_clock = clock;
  assign RetimeWrapper_72_reset = reset;
  assign _T_2952 = RetimeWrapper_72_io_out;
  assign RetimeWrapper_73_io_flow = 1'h1;
  assign RetimeWrapper_73_io_in = x3300_sm_io_output_rst_en;
  assign RetimeWrapper_73_clock = clock;
  assign RetimeWrapper_73_reset = reset;
  assign _T_2961 = RetimeWrapper_73_io_out;
  assign RetimeWrapper_74_io_flow = 1'h1;
  assign RetimeWrapper_74_io_in = x3300_sm_io_output_stageEnable_1;
  assign RetimeWrapper_74_clock = clock;
  assign RetimeWrapper_74_reset = reset;
  assign _T_2967 = RetimeWrapper_74_io_out;
  assign RetimeWrapper_75_io_flow = 1'h1;
  assign RetimeWrapper_75_io_in = _T_2970;
  assign RetimeWrapper_75_clock = clock;
  assign RetimeWrapper_75_reset = reset;
  assign _T_2974 = RetimeWrapper_75_io_out;
  assign RetimeWrapper_76_io_flow = 1'h1;
  assign RetimeWrapper_76_io_in = x3300_sm_io_output_rst_en;
  assign RetimeWrapper_76_clock = clock;
  assign RetimeWrapper_76_reset = reset;
  assign _T_2981 = RetimeWrapper_76_io_out;
  assign RetimeWrapper_77_io_flow = _T_2986;
  assign RetimeWrapper_77_io_in = _T_3002;
  assign RetimeWrapper_77_clock = clock;
  assign RetimeWrapper_77_reset = reset;
  assign _T_3007 = RetimeWrapper_77_io_out;
  assign RetimeWrapper_78_io_flow = _T_2986;
  assign RetimeWrapper_78_io_in = x3237_ctr_trivial;
  assign RetimeWrapper_78_clock = clock;
  assign RetimeWrapper_78_reset = reset;
  assign _T_3016 = RetimeWrapper_78_io_out;
  assign RetimeWrapper_79_io_flow = 1'h1;
  assign RetimeWrapper_79_io_in = x3237_ctr_trivial;
  assign RetimeWrapper_79_clock = clock;
  assign RetimeWrapper_79_reset = reset;
  assign _T_3048 = RetimeWrapper_79_io_out;
  assign RetimeWrapper_80_io_flow = 1'h1;
  assign RetimeWrapper_80_io_in = x3236_sm_io_output_stageEnable_0;
  assign RetimeWrapper_80_clock = clock;
  assign RetimeWrapper_80_reset = reset;
  assign _T_3056 = RetimeWrapper_80_io_out;
  assign RetimeWrapper_81_io_flow = 1'h1;
  assign RetimeWrapper_81_io_in = _T_3059;
  assign RetimeWrapper_81_clock = clock;
  assign RetimeWrapper_81_reset = reset;
  assign _T_3063 = RetimeWrapper_81_io_out;
  assign RetimeWrapper_82_io_flow = 1'h1;
  assign RetimeWrapper_82_io_in = _T_3067;
  assign RetimeWrapper_82_clock = clock;
  assign RetimeWrapper_82_reset = reset;
  assign _T_3071 = RetimeWrapper_82_io_out;
  assign RetimeWrapper_83_io_flow = 1'h1;
  assign RetimeWrapper_83_io_in = x3236_sm_io_output_rst_en;
  assign RetimeWrapper_83_clock = clock;
  assign RetimeWrapper_83_reset = reset;
  assign _T_3080 = RetimeWrapper_83_io_out;
  assign RetimeWrapper_84_io_flow = 1'h1;
  assign RetimeWrapper_84_io_in = x3236_sm_io_output_stageEnable_1;
  assign RetimeWrapper_84_clock = clock;
  assign RetimeWrapper_84_reset = reset;
  assign _T_3086 = RetimeWrapper_84_io_out;
  assign RetimeWrapper_85_io_flow = 1'h1;
  assign RetimeWrapper_85_io_in = _T_3089;
  assign RetimeWrapper_85_clock = clock;
  assign RetimeWrapper_85_reset = reset;
  assign _T_3093 = RetimeWrapper_85_io_out;
  assign RetimeWrapper_86_io_flow = 1'h1;
  assign RetimeWrapper_86_io_in = x3236_sm_io_output_rst_en;
  assign RetimeWrapper_86_clock = clock;
  assign RetimeWrapper_86_reset = reset;
  assign RetimeWrapper_87_io_flow = 1'h1;
  assign RetimeWrapper_87_io_in = _T_3121;
  assign RetimeWrapper_87_clock = clock;
  assign RetimeWrapper_87_reset = reset;
  assign _T_3125 = RetimeWrapper_87_io_out;
  assign RetimeWrapper_88_io_flow = 1'h1;
  assign RetimeWrapper_88_io_in = x3236_ctr_trivial;
  assign RetimeWrapper_88_clock = clock;
  assign RetimeWrapper_88_reset = reset;
  assign _T_3133 = RetimeWrapper_88_io_out;
  assign RetimeWrapper_89_io_flow = 1'h1;
  assign RetimeWrapper_89_io_in = x3235_done;
  assign RetimeWrapper_89_clock = clock;
  assign RetimeWrapper_89_reset = reset;
  assign _T_3419 = RetimeWrapper_89_io_out;
  assign RetimeWrapper_90_io_flow = 1'h1;
  assign RetimeWrapper_90_io_in = x3223_done;
  assign RetimeWrapper_90_clock = clock;
  assign RetimeWrapper_90_reset = reset;
  assign _T_3425 = RetimeWrapper_90_io_out;
  assign _T_3504_number = _T_3514;
  assign _T_3506_number = _T_3525;
  assign _T_3514 = b1270_number;
  assign _T_3525 = x3221_number;
  assign RetimeWrapper_91_io_flow = 1'h1;
  assign RetimeWrapper_91_io_in = x3236_ctr_trivial;
  assign RetimeWrapper_91_clock = clock;
  assign RetimeWrapper_91_reset = reset;
  assign _T_3565 = RetimeWrapper_91_io_out;
  assign _T_3569_number = _T_3579;
  assign _T_3579 = x3221_number;
  assign RetimeWrapper_92_io_flow = 1'h1;
  assign RetimeWrapper_92_io_in = x3428_ctr_trivial;
  assign RetimeWrapper_92_clock = clock;
  assign RetimeWrapper_92_reset = reset;
  assign _T_3609 = RetimeWrapper_92_io_out;
  assign RetimeWrapper_93_io_flow = 1'h1;
  assign RetimeWrapper_93_io_in = x3364_sm_io_output_stageEnable_0;
  assign RetimeWrapper_93_clock = clock;
  assign RetimeWrapper_93_reset = reset;
  assign _T_3617 = RetimeWrapper_93_io_out;
  assign RetimeWrapper_94_io_flow = 1'h1;
  assign RetimeWrapper_94_io_in = _T_3620;
  assign RetimeWrapper_94_clock = clock;
  assign RetimeWrapper_94_reset = reset;
  assign _T_3624 = RetimeWrapper_94_io_out;
  assign RetimeWrapper_95_io_flow = 1'h1;
  assign RetimeWrapper_95_io_in = _T_3629;
  assign RetimeWrapper_95_clock = clock;
  assign RetimeWrapper_95_reset = reset;
  assign _T_3633 = RetimeWrapper_95_io_out;
  assign RetimeWrapper_96_io_flow = 1'h1;
  assign RetimeWrapper_96_io_in = x3364_sm_io_output_rst_en;
  assign RetimeWrapper_96_clock = clock;
  assign RetimeWrapper_96_reset = reset;
  assign _T_3642 = RetimeWrapper_96_io_out;
  assign RetimeWrapper_97_io_flow = 1'h1;
  assign RetimeWrapper_97_io_in = x3364_sm_io_output_stageEnable_1;
  assign RetimeWrapper_97_clock = clock;
  assign RetimeWrapper_97_reset = reset;
  assign _T_3648 = RetimeWrapper_97_io_out;
  assign RetimeWrapper_98_io_flow = 1'h1;
  assign RetimeWrapper_98_io_in = _T_3651;
  assign RetimeWrapper_98_clock = clock;
  assign RetimeWrapper_98_reset = reset;
  assign _T_3655 = RetimeWrapper_98_io_out;
  assign RetimeWrapper_99_io_flow = 1'h1;
  assign RetimeWrapper_99_io_in = x3364_sm_io_output_rst_en;
  assign RetimeWrapper_99_clock = clock;
  assign RetimeWrapper_99_reset = reset;
  assign _T_3662 = RetimeWrapper_99_io_out;
  assign RetimeWrapper_100_io_flow = 1'h1;
  assign RetimeWrapper_100_io_in = x3428_ctr_trivial;
  assign RetimeWrapper_100_clock = clock;
  assign RetimeWrapper_100_reset = reset;
  assign _T_3678 = RetimeWrapper_100_io_out;
  assign RetimeWrapper_101_io_flow = 1'h1;
  assign RetimeWrapper_101_io_in = x3427_sm_io_output_stageEnable_0;
  assign RetimeWrapper_101_clock = clock;
  assign RetimeWrapper_101_reset = reset;
  assign _T_3686 = RetimeWrapper_101_io_out;
  assign RetimeWrapper_102_io_flow = 1'h1;
  assign RetimeWrapper_102_io_in = _T_3689;
  assign RetimeWrapper_102_clock = clock;
  assign RetimeWrapper_102_reset = reset;
  assign _T_3693 = RetimeWrapper_102_io_out;
  assign RetimeWrapper_103_io_flow = 1'h1;
  assign RetimeWrapper_103_io_in = _T_3698;
  assign RetimeWrapper_103_clock = clock;
  assign RetimeWrapper_103_reset = reset;
  assign _T_3702 = RetimeWrapper_103_io_out;
  assign RetimeWrapper_104_io_flow = 1'h1;
  assign RetimeWrapper_104_io_in = x3427_sm_io_output_rst_en;
  assign RetimeWrapper_104_clock = clock;
  assign RetimeWrapper_104_reset = reset;
  assign _T_3711 = RetimeWrapper_104_io_out;
  assign RetimeWrapper_105_io_flow = 1'h1;
  assign RetimeWrapper_105_io_in = x3427_sm_io_output_stageEnable_1;
  assign RetimeWrapper_105_clock = clock;
  assign RetimeWrapper_105_reset = reset;
  assign _T_3717 = RetimeWrapper_105_io_out;
  assign RetimeWrapper_106_io_flow = 1'h1;
  assign RetimeWrapper_106_io_in = _T_3720;
  assign RetimeWrapper_106_clock = clock;
  assign RetimeWrapper_106_reset = reset;
  assign _T_3724 = RetimeWrapper_106_io_out;
  assign RetimeWrapper_107_io_flow = 1'h1;
  assign RetimeWrapper_107_io_in = x3427_sm_io_output_rst_en;
  assign RetimeWrapper_107_clock = clock;
  assign RetimeWrapper_107_reset = reset;
  assign _T_3731 = RetimeWrapper_107_io_out;
  assign RetimeWrapper_108_io_flow = _T_3736;
  assign RetimeWrapper_108_io_in = _T_3752;
  assign RetimeWrapper_108_clock = clock;
  assign RetimeWrapper_108_reset = reset;
  assign _T_3757 = RetimeWrapper_108_io_out;
  assign RetimeWrapper_109_io_flow = _T_3736;
  assign RetimeWrapper_109_io_in = x3427_ctr_trivial;
  assign RetimeWrapper_109_clock = clock;
  assign RetimeWrapper_109_reset = reset;
  assign _T_3766 = RetimeWrapper_109_io_out;
  assign RetimeWrapper_110_io_flow = 1'h1;
  assign RetimeWrapper_110_io_in = x3427_ctr_trivial;
  assign RetimeWrapper_110_clock = clock;
  assign RetimeWrapper_110_reset = reset;
  assign _T_3798 = RetimeWrapper_110_io_out;
  assign RetimeWrapper_111_io_flow = 1'h1;
  assign RetimeWrapper_111_io_in = x3426_sm_io_output_stageEnable_0;
  assign RetimeWrapper_111_clock = clock;
  assign RetimeWrapper_111_reset = reset;
  assign _T_3806 = RetimeWrapper_111_io_out;
  assign RetimeWrapper_112_io_flow = 1'h1;
  assign RetimeWrapper_112_io_in = _T_3809;
  assign RetimeWrapper_112_clock = clock;
  assign RetimeWrapper_112_reset = reset;
  assign _T_3813 = RetimeWrapper_112_io_out;
  assign RetimeWrapper_113_io_flow = 1'h1;
  assign RetimeWrapper_113_io_in = _T_3817;
  assign RetimeWrapper_113_clock = clock;
  assign RetimeWrapper_113_reset = reset;
  assign _T_3821 = RetimeWrapper_113_io_out;
  assign RetimeWrapper_114_io_flow = 1'h1;
  assign RetimeWrapper_114_io_in = x3426_sm_io_output_rst_en;
  assign RetimeWrapper_114_clock = clock;
  assign RetimeWrapper_114_reset = reset;
  assign _T_3830 = RetimeWrapper_114_io_out;
  assign RetimeWrapper_115_io_flow = 1'h1;
  assign RetimeWrapper_115_io_in = x3426_sm_io_output_stageEnable_1;
  assign RetimeWrapper_115_clock = clock;
  assign RetimeWrapper_115_reset = reset;
  assign _T_3836 = RetimeWrapper_115_io_out;
  assign RetimeWrapper_116_io_flow = 1'h1;
  assign RetimeWrapper_116_io_in = _T_3839;
  assign RetimeWrapper_116_clock = clock;
  assign RetimeWrapper_116_reset = reset;
  assign _T_3843 = RetimeWrapper_116_io_out;
  assign RetimeWrapper_117_io_flow = 1'h1;
  assign RetimeWrapper_117_io_in = x3426_sm_io_output_rst_en;
  assign RetimeWrapper_117_clock = clock;
  assign RetimeWrapper_117_reset = reset;
  assign _T_3855_number = _T_3865;
  assign _T_3857_number = b1202_chain_read_1;
  assign _T_3865 = _T_3857_number;
  assign _T_3870_number = _T_3871[31:0];
  assign _T_3873_number = _T_3874[31:0];
  assign _T_3876_number = _T_3909;
  assign _T_3878_number = _T_3888;
  assign _T_3880_number = _T_3901;
  assign _T_3888 = _T_3893;
  assign _T_3901 = _T_3906;
  assign _T_3911_number = _T_3925;
  assign _T_3925 = _T_3929;
  assign _T_3931_number = _T_3963;
  assign _T_3933_number = _T_3943;
  assign _T_3935_number = _T_3956;
  assign _T_3943 = _T_3893;
  assign _T_3956 = _T_3961;
  assign _T_3965_number = _T_3979;
  assign _T_3979 = _T_3983;
  assign _T_3989_number = _T_3999;
  assign _T_3999 = x3189_number;
  assign _T_4020_number = _T_4053;
  assign _T_4024_number = _T_4045;
  assign _T_4045 = _T_4050;
  assign _T_4055_number = _T_4069;
  assign _T_4069 = _T_4073;
  assign _T_4080_number = _T_4087;
  assign _T_4089_number = _T_4096;
  assign _T_4098_number = _T_4130;
  assign _T_4100_number = _T_4110;
  assign _T_4102_number = _T_4123;
  assign _T_4110 = _T_4115;
  assign _T_4123 = _T_4128;
  assign _T_4132_number = _T_4146;
  assign _T_4146 = _T_4150;
  assign _T_4152_number = _T_4184;
  assign _T_4154_number = _T_4164;
  assign _T_4156_number = _T_4177;
  assign _T_4164 = _T_4128;
  assign _T_4177 = _T_4115;
  assign _T_4186_number = _T_4200;
  assign _T_4200 = _T_4204;
  assign _T_4206_number = _T_4238;
  assign _T_4208_number = _T_4218;
  assign _T_4210_number = _T_4231;
  assign _T_4218 = _T_4223;
  assign _T_4231 = _T_4236;
  assign _T_4240_number = _T_4254;
  assign _T_4254 = _T_4258;
  assign _T_4260_number = _T_4292;
  assign _T_4262_number = _T_4272;
  assign _T_4264_number = _T_4285;
  assign _T_4272 = _T_3961;
  assign _T_4285 = _T_3906;
  assign _T_4294_number = _T_4308;
  assign _T_4308 = _T_4312;
  assign _T_4314_number = _T_4346;
  assign _T_4316_number = _T_4326;
  assign _T_4318_number = _T_4339;
  assign _T_4326 = _T_4331;
  assign _T_4339 = _T_4344;
  assign _T_4348_number = _T_4362;
  assign _T_4362 = _T_4366;
  assign _T_4374 = _T_4383;
  assign _T_4385_number = _T_4395;
  assign _T_4387_number = io_argIns_1;
  assign _T_4395 = _T_4387_number;
  assign _T_4400_number = _T_4432;
  assign _T_4402_number = _T_4412;
  assign _T_4404_number = _T_4425;
  assign _T_4412 = _T_4417;
  assign _T_4425 = _T_4430;
  assign _T_4434_number = _T_4448;
  assign _T_4448 = _T_4452;
  assign _T_4460 = x3202_number;
  assign _T_4485_0 = x3206;
  assign _T_4499_0 = _T_4473;
  assign RetimeWrapper_118_io_flow = _T_4505;
  assign RetimeWrapper_118_io_in = _T_4521;
  assign RetimeWrapper_118_clock = clock;
  assign RetimeWrapper_118_reset = reset;
  assign _T_4526 = RetimeWrapper_118_io_out;
  assign RetimeWrapper_119_io_flow = _T_4505;
  assign RetimeWrapper_119_io_in = x3300_ctr_trivial;
  assign RetimeWrapper_119_clock = clock;
  assign RetimeWrapper_119_reset = reset;
  assign _T_4535 = RetimeWrapper_119_io_out;
  assign RetimeWrapper_120_io_flow = 1'h1;
  assign RetimeWrapper_120_io_in = x3300_ctr_trivial;
  assign RetimeWrapper_120_clock = clock;
  assign RetimeWrapper_120_reset = reset;
  assign _T_4567 = RetimeWrapper_120_io_out;
  assign RetimeWrapper_121_io_flow = 1'h1;
  assign RetimeWrapper_121_io_in = x3299_sm_io_output_stageEnable_0;
  assign RetimeWrapper_121_clock = clock;
  assign RetimeWrapper_121_reset = reset;
  assign _T_4575 = RetimeWrapper_121_io_out;
  assign RetimeWrapper_122_io_flow = 1'h1;
  assign RetimeWrapper_122_io_in = _T_4578;
  assign RetimeWrapper_122_clock = clock;
  assign RetimeWrapper_122_reset = reset;
  assign _T_4582 = RetimeWrapper_122_io_out;
  assign RetimeWrapper_123_io_flow = 1'h1;
  assign RetimeWrapper_123_io_in = _T_4586;
  assign RetimeWrapper_123_clock = clock;
  assign RetimeWrapper_123_reset = reset;
  assign _T_4590 = RetimeWrapper_123_io_out;
  assign RetimeWrapper_124_io_flow = 1'h1;
  assign RetimeWrapper_124_io_in = x3299_sm_io_output_rst_en;
  assign RetimeWrapper_124_clock = clock;
  assign RetimeWrapper_124_reset = reset;
  assign _T_4599 = RetimeWrapper_124_io_out;
  assign RetimeWrapper_125_io_flow = 1'h1;
  assign RetimeWrapper_125_io_in = x3299_sm_io_output_stageEnable_1;
  assign RetimeWrapper_125_clock = clock;
  assign RetimeWrapper_125_reset = reset;
  assign _T_4605 = RetimeWrapper_125_io_out;
  assign RetimeWrapper_126_io_flow = 1'h1;
  assign RetimeWrapper_126_io_in = _T_4608;
  assign RetimeWrapper_126_clock = clock;
  assign RetimeWrapper_126_reset = reset;
  assign _T_4612 = RetimeWrapper_126_io_out;
  assign RetimeWrapper_127_io_flow = 1'h1;
  assign RetimeWrapper_127_io_in = x3299_sm_io_output_rst_en;
  assign RetimeWrapper_127_clock = clock;
  assign RetimeWrapper_127_reset = reset;
  assign RetimeWrapper_128_io_flow = 1'h1;
  assign RetimeWrapper_128_io_in = _T_4640;
  assign RetimeWrapper_128_clock = clock;
  assign RetimeWrapper_128_reset = reset;
  assign _T_4644 = RetimeWrapper_128_io_out;
  assign RetimeWrapper_129_io_flow = 1'h1;
  assign RetimeWrapper_129_io_in = x3299_ctr_trivial;
  assign RetimeWrapper_129_clock = clock;
  assign RetimeWrapper_129_reset = reset;
  assign _T_4652 = RetimeWrapper_129_io_out;
  assign RetimeWrapper_130_io_flow = 1'h1;
  assign RetimeWrapper_130_io_in = x3298_done;
  assign RetimeWrapper_130_clock = clock;
  assign RetimeWrapper_130_reset = reset;
  assign _T_4938 = RetimeWrapper_130_io_out;
  assign RetimeWrapper_131_io_flow = 1'h1;
  assign RetimeWrapper_131_io_in = x3286_done;
  assign RetimeWrapper_131_clock = clock;
  assign RetimeWrapper_131_reset = reset;
  assign _T_4944 = RetimeWrapper_131_io_out;
  assign _T_5023_number = _T_5033;
  assign _T_5025_number = _T_5044;
  assign _T_5033 = b1331_number;
  assign _T_5044 = x3284_number;
  assign RetimeWrapper_132_io_flow = 1'h1;
  assign RetimeWrapper_132_io_in = x3299_ctr_trivial;
  assign RetimeWrapper_132_clock = clock;
  assign RetimeWrapper_132_reset = reset;
  assign _T_5084 = RetimeWrapper_132_io_out;
  assign _T_5088_number = _T_5098;
  assign _T_5098 = x3284_number;
  assign RetimeWrapper_133_io_flow = 1'h1;
  assign RetimeWrapper_133_io_in = x3433_done;
  assign RetimeWrapper_133_clock = clock;
  assign RetimeWrapper_133_reset = reset;
  assign _T_5407 = RetimeWrapper_133_io_out;
  assign _T_5491_number = _T_5501;
  assign _T_5493_number = _T_5512;
  assign _T_5501 = b1479_number;
  assign _T_5512 = x3431_number;
  assign _T_5621_number = _T_5631;
  assign _T_5623_number = _T_5642;
  assign _T_5631 = b1480_number;
  assign _T_5642 = x3431_number;
  assign _T_5751_number = _T_5761;
  assign _T_5753_number = _T_5772;
  assign _T_5761 = b1481_number;
  assign _T_5772 = x3431_number;
  assign _T_5881_number = _T_5891;
  assign _T_5883_number = _T_5902;
  assign _T_5891 = b1482_number;
  assign _T_5902 = x3431_number;
  assign RetimeWrapper_134_io_flow = 1'h1;
  assign RetimeWrapper_134_io_in = x3503_ctr_trivial;
  assign RetimeWrapper_134_clock = clock;
  assign RetimeWrapper_134_reset = reset;
  assign _T_5942 = RetimeWrapper_134_io_out;
  assign _T_5946_number = _T_5956;
  assign _T_5956 = x3431_number;
  assign RetimeWrapper_135_io_flow = 1'h1;
  assign RetimeWrapper_135_io_in = x3469_done;
  assign RetimeWrapper_135_clock = clock;
  assign RetimeWrapper_135_reset = reset;
  assign _T_6265 = RetimeWrapper_135_io_out;
  assign _T_6349_number = _T_6359;
  assign _T_6351_number = _T_6370;
  assign _T_6359 = b1520_number;
  assign _T_6370 = x3467_number;
  assign _T_6479_number = _T_6489;
  assign _T_6481_number = _T_6500;
  assign _T_6489 = b1521_number;
  assign _T_6500 = x3467_number;
  assign _T_6609_number = _T_6619;
  assign _T_6611_number = _T_6630;
  assign _T_6619 = b1522_number;
  assign _T_6630 = x3467_number;
  assign _T_6739_number = _T_6749;
  assign _T_6741_number = _T_6760;
  assign _T_6749 = b1523_number;
  assign _T_6760 = x3467_number;
  assign RetimeWrapper_136_io_flow = 1'h1;
  assign RetimeWrapper_136_io_in = x3503_ctr_trivial;
  assign RetimeWrapper_136_clock = clock;
  assign RetimeWrapper_136_reset = reset;
  assign _T_6800 = RetimeWrapper_136_io_out;
  assign _T_6804_number = _T_6814;
  assign _T_6814 = x3467_number;
  assign _T_6832_number = _T_6864;
  assign _T_6834_number = _T_6849;
  assign _T_6836_number = _T_6862;
  assign _T_6840 = _T_6845;
  assign _T_6842 = _T_6840;
  assign _T_6844 = _T_6848;
  assign _T_6853 = _T_6858;
  assign _T_6855 = _T_6853;
  assign _T_6857 = _T_6861;
  assign _T_6866_number = _T_6884;
  assign _T_6876 = _T_6881;
  assign _T_6878 = _T_6876;
  assign _T_6880 = _T_6883;
  assign _T_6894_number = _T_6904;
  assign _T_6896_number = b1202_chain_read_4;
  assign _T_6904 = _T_6896_number;
  assign _T_6909_number = _T_6919;
  assign _T_6919 = _T_6894_number;
  assign _T_6936_number = _T_6968;
  assign _T_6938_number = _T_6953;
  assign _T_6944 = _T_6949;
  assign _T_6946 = _T_6944;
  assign _T_6948 = _T_6952;
  assign _T_6970_number = _T_6988;
  assign _T_6980 = _T_6985;
  assign _T_6982 = _T_6980;
  assign _T_6984 = _T_6987;
  assign RetimeWrapper_137_io_flow = 1'h1;
  assign RetimeWrapper_137_io_in = x3152_wren;
  assign RetimeWrapper_137_clock = clock;
  assign RetimeWrapper_137_reset = reset;
  assign _T_6995 = RetimeWrapper_137_io_out;
  assign RetimeWrapper_138_io_flow = 1'h1;
  assign RetimeWrapper_138_io_in = reset;
  assign RetimeWrapper_138_clock = clock;
  assign RetimeWrapper_138_reset = reset;
  assign _T_7002 = RetimeWrapper_138_io_out;
  assign _T_7020_number = _T_7030;
  assign _T_7022_number = b1203_chain_read_1;
  assign _T_7030 = _T_7022_number;
  assign _T_7035_number = _T_7036[31:0];
  assign _T_7038_number = _T_7039[31:0];
  assign _T_7041_number = _T_7074;
  assign _T_7043_number = _T_7053;
  assign _T_7045_number = _T_7066;
  assign _T_7053 = _T_7058;
  assign _T_7066 = _T_7071;
  assign _T_7076_number = _T_7090;
  assign _T_7090 = _T_7094;
  assign _T_7096_number = _T_7128;
  assign _T_7098_number = _T_7108;
  assign _T_7100_number = _T_7121;
  assign _T_7108 = _T_7058;
  assign _T_7121 = _T_7126;
  assign _T_7130_number = _T_7144;
  assign _T_7144 = _T_7148;
  assign _T_7154_number = _T_7164;
  assign _T_7164 = x3252_number;
  assign _T_7185_number = _T_7218;
  assign _T_7189_number = _T_7210;
  assign _T_7210 = _T_7215;
  assign _T_7220_number = _T_7234;
  assign _T_7234 = _T_7238;
  assign _T_7245_number = _T_7252;
  assign _T_7254_number = _T_7261;
  assign _T_7263_number = _T_7295;
  assign _T_7265_number = _T_7275;
  assign _T_7267_number = _T_7288;
  assign _T_7275 = _T_7280;
  assign _T_7288 = _T_7293;
  assign _T_7297_number = _T_7311;
  assign _T_7311 = _T_7315;
  assign _T_7317_number = _T_7349;
  assign _T_7319_number = _T_7329;
  assign _T_7321_number = _T_7342;
  assign _T_7329 = _T_7293;
  assign _T_7342 = _T_7280;
  assign _T_7351_number = _T_7365;
  assign _T_7365 = _T_7369;
  assign _T_7371_number = _T_7403;
  assign _T_7373_number = _T_7383;
  assign _T_7375_number = _T_7396;
  assign _T_7383 = _T_7388;
  assign _T_7396 = _T_7401;
  assign _T_7405_number = _T_7419;
  assign _T_7419 = _T_7423;
  assign _T_7425_number = _T_7457;
  assign _T_7427_number = _T_7437;
  assign _T_7429_number = _T_7450;
  assign _T_7437 = _T_7126;
  assign _T_7450 = _T_7071;
  assign _T_7459_number = _T_7473;
  assign _T_7473 = _T_7477;
  assign _T_7479_number = _T_7511;
  assign _T_7481_number = _T_7491;
  assign _T_7483_number = _T_7504;
  assign _T_7491 = _T_7496;
  assign _T_7504 = _T_7509;
  assign _T_7513_number = _T_7527;
  assign _T_7527 = _T_7531;
  assign _T_7539 = _T_7548;
  assign _T_7550_number = _T_7560;
  assign _T_7552_number = io_argIns_1;
  assign _T_7560 = _T_7552_number;
  assign _T_7565_number = _T_7597;
  assign _T_7567_number = _T_7577;
  assign _T_7569_number = _T_7590;
  assign _T_7577 = _T_7582;
  assign _T_7590 = _T_7595;
  assign _T_7599_number = _T_7613;
  assign _T_7613 = _T_7617;
  assign _T_7625 = x3265_number;
  assign _T_7650_0 = x3269;
  assign _T_7664_0 = _T_7638;
  assign _T_7669_number = _T_7679;
  assign _T_7671_number = b1203_chain_read_2;
  assign _T_7679 = _T_7671_number;
  assign _T_7684_number = _T_7685[31:0];
  assign _T_7687_number = _T_7688[31:0];
  assign _T_7690_number = _T_7723;
  assign _T_7692_number = _T_7702;
  assign _T_7694_number = _T_7715;
  assign _T_7702 = _T_7707;
  assign _T_7715 = _T_7720;
  assign _T_7725_number = _T_7739;
  assign _T_7739 = _T_7743;
  assign _T_7745_number = _T_7777;
  assign _T_7747_number = _T_7757;
  assign _T_7749_number = _T_7770;
  assign _T_7757 = _T_7707;
  assign _T_7770 = _T_7775;
  assign _T_7779_number = _T_7793;
  assign _T_7793 = _T_7797;
  assign _T_7803_number = _T_7813;
  assign _T_7813 = x3379_number;
  assign _T_7834_number = _T_7867;
  assign _T_7838_number = _T_7859;
  assign _T_7859 = _T_7864;
  assign _T_7869_number = _T_7883;
  assign _T_7883 = _T_7887;
  assign _T_7894_number = _T_7901;
  assign _T_7903_number = _T_7910;
  assign _T_7912_number = _T_7944;
  assign _T_7914_number = _T_7924;
  assign _T_7916_number = _T_7937;
  assign _T_7924 = _T_7929;
  assign _T_7937 = _T_7942;
  assign _T_7946_number = _T_7960;
  assign _T_7960 = _T_7964;
  assign _T_7966_number = _T_7998;
  assign _T_7968_number = _T_7978;
  assign _T_7970_number = _T_7991;
  assign _T_7978 = _T_7942;
  assign _T_7991 = _T_7929;
  assign _T_8000_number = _T_8014;
  assign _T_8014 = _T_8018;
  assign _T_8020_number = _T_8052;
  assign _T_8022_number = _T_8032;
  assign _T_8024_number = _T_8045;
  assign _T_8032 = _T_8037;
  assign _T_8045 = _T_8050;
  assign _T_8054_number = _T_8068;
  assign _T_8068 = _T_8072;
  assign _T_8074_number = _T_8106;
  assign _T_8076_number = _T_8086;
  assign _T_8078_number = _T_8099;
  assign _T_8086 = _T_7775;
  assign _T_8099 = _T_7720;
  assign _T_8108_number = _T_8122;
  assign _T_8122 = _T_8126;
  assign _T_8128_number = _T_8160;
  assign _T_8130_number = _T_8140;
  assign _T_8132_number = _T_8153;
  assign _T_8140 = _T_8145;
  assign _T_8153 = _T_8158;
  assign _T_8162_number = _T_8176;
  assign _T_8176 = _T_8180;
  assign _T_8188 = _T_8197;
  assign _T_8199_number = _T_8209;
  assign _T_8201_number = io_argIns_2;
  assign _T_8209 = _T_8201_number;
  assign _T_8214_number = _T_8246;
  assign _T_8216_number = _T_8226;
  assign _T_8218_number = _T_8239;
  assign _T_8226 = _T_8231;
  assign _T_8239 = _T_8244;
  assign _T_8248_number = _T_8262;
  assign _T_8262 = _T_8266;
  assign _T_8274 = x3392_number;
  assign _T_8299_0 = x3396;
  assign _T_8313_0 = _T_8287;
  assign RetimeWrapper_139_io_flow = 1'h1;
  assign RetimeWrapper_139_io_in = _T_8345;
  assign RetimeWrapper_139_clock = clock;
  assign RetimeWrapper_139_reset = reset;
  assign _T_8349 = RetimeWrapper_139_io_out;
  assign RetimeWrapper_140_io_flow = 1'h1;
  assign RetimeWrapper_140_io_in = x3174_ctr_trivial;
  assign RetimeWrapper_140_clock = clock;
  assign RetimeWrapper_140_reset = reset;
  assign _T_8357 = RetimeWrapper_140_io_out;
  assign RetimeWrapper_141_io_flow = 1'h1;
  assign RetimeWrapper_141_io_in = _T_8391;
  assign RetimeWrapper_141_clock = clock;
  assign RetimeWrapper_141_reset = reset;
  assign _T_8395 = RetimeWrapper_141_io_out;
  assign RetimeWrapper_142_io_flow = 1'h1;
  assign RetimeWrapper_142_io_in = x3174_ctr_trivial;
  assign RetimeWrapper_142_clock = clock;
  assign RetimeWrapper_142_reset = reset;
  assign _T_8403 = RetimeWrapper_142_io_out;
  assign _T_8410_number = _T_8443;
  assign _T_8412_number = _T_8422;
  assign _T_8414_number = _T_8435;
  assign _T_8422 = _T_8427;
  assign _T_8435 = _T_8440;
  assign _T_8445_number = _T_8459;
  assign _T_8459 = _T_8463;
  assign _T_8471_number = _T_8490;
  assign _T_8490 = x3169_number;
  assign RetimeWrapper_143_io_flow = 1'h1;
  assign RetimeWrapper_143_io_in = reset;
  assign RetimeWrapper_143_clock = clock;
  assign RetimeWrapper_143_reset = reset;
  assign _T_8564 = RetimeWrapper_143_io_out;
  assign RetimeWrapper_144_io_flow = 1'h1;
  assign RetimeWrapper_144_io_in = x3174_done;
  assign RetimeWrapper_144_clock = clock;
  assign RetimeWrapper_144_reset = reset;
  assign _T_8571 = RetimeWrapper_144_io_out;
  assign RetimeWrapper_145_io_flow = 1'h1;
  assign RetimeWrapper_145_io_in = x3301_done;
  assign RetimeWrapper_145_clock = clock;
  assign RetimeWrapper_145_reset = reset;
  assign _T_8577 = RetimeWrapper_145_io_out;
  assign RetimeWrapper_146_io_flow = 1'h1;
  assign RetimeWrapper_146_io_in = x3428_done;
  assign RetimeWrapper_146_clock = clock;
  assign RetimeWrapper_146_reset = reset;
  assign _T_8583 = RetimeWrapper_146_io_out;
  assign RetimeWrapper_147_io_flow = 1'h1;
  assign RetimeWrapper_147_io_in = x3503_done;
  assign RetimeWrapper_147_clock = clock;
  assign RetimeWrapper_147_reset = reset;
  assign _T_8589 = RetimeWrapper_147_io_out;
  assign RetimeWrapper_148_io_flow = 1'h1;
  assign RetimeWrapper_148_io_in = x3514_done;
  assign RetimeWrapper_148_clock = clock;
  assign RetimeWrapper_148_reset = reset;
  assign _T_8595 = RetimeWrapper_148_io_out;
  assign RetimeWrapper_149_io_flow = 1'h1;
  assign RetimeWrapper_149_io_in = x3174_done;
  assign RetimeWrapper_149_clock = clock;
  assign RetimeWrapper_149_reset = reset;
  assign _T_8601 = RetimeWrapper_149_io_out;
  assign RetimeWrapper_150_io_flow = 1'h1;
  assign RetimeWrapper_150_io_in = x3301_done;
  assign RetimeWrapper_150_clock = clock;
  assign RetimeWrapper_150_reset = reset;
  assign _T_8607 = RetimeWrapper_150_io_out;
  assign RetimeWrapper_151_io_flow = 1'h1;
  assign RetimeWrapper_151_io_in = x3428_done;
  assign RetimeWrapper_151_clock = clock;
  assign RetimeWrapper_151_reset = reset;
  assign _T_8613 = RetimeWrapper_151_io_out;
  assign RetimeWrapper_152_io_flow = 1'h1;
  assign RetimeWrapper_152_io_in = x3503_done;
  assign RetimeWrapper_152_clock = clock;
  assign RetimeWrapper_152_reset = reset;
  assign _T_8619 = RetimeWrapper_152_io_out;
  assign RetimeWrapper_153_io_flow = 1'h1;
  assign RetimeWrapper_153_io_in = x3514_done;
  assign RetimeWrapper_153_clock = clock;
  assign RetimeWrapper_153_reset = reset;
  assign _T_8625 = RetimeWrapper_153_io_out;
  assign RetimeWrapper_154_io_flow = 1'h1;
  assign RetimeWrapper_154_io_in = x3174_done;
  assign RetimeWrapper_154_clock = clock;
  assign RetimeWrapper_154_reset = reset;
  assign _T_8661 = RetimeWrapper_154_io_out;
  assign RetimeWrapper_155_io_flow = 1'h1;
  assign RetimeWrapper_155_io_in = x3301_done;
  assign RetimeWrapper_155_clock = clock;
  assign RetimeWrapper_155_reset = reset;
  assign _T_8667 = RetimeWrapper_155_io_out;
  assign RetimeWrapper_156_io_flow = 1'h1;
  assign RetimeWrapper_156_io_in = x3428_done;
  assign RetimeWrapper_156_clock = clock;
  assign RetimeWrapper_156_reset = reset;
  assign _T_8673 = RetimeWrapper_156_io_out;
  assign RetimeWrapper_157_io_flow = 1'h1;
  assign RetimeWrapper_157_io_in = x3503_done;
  assign RetimeWrapper_157_clock = clock;
  assign RetimeWrapper_157_reset = reset;
  assign _T_8679 = RetimeWrapper_157_io_out;
  assign RetimeWrapper_158_io_flow = 1'h1;
  assign RetimeWrapper_158_io_in = x3174_done;
  assign RetimeWrapper_158_clock = clock;
  assign RetimeWrapper_158_reset = reset;
  assign _T_8685 = RetimeWrapper_158_io_out;
  assign RetimeWrapper_159_io_flow = 1'h1;
  assign RetimeWrapper_159_io_in = x3301_done;
  assign RetimeWrapper_159_clock = clock;
  assign RetimeWrapper_159_reset = reset;
  assign _T_8691 = RetimeWrapper_159_io_out;
  assign RetimeWrapper_160_io_flow = 1'h1;
  assign RetimeWrapper_160_io_in = x3428_done;
  assign RetimeWrapper_160_clock = clock;
  assign RetimeWrapper_160_reset = reset;
  assign _T_8697 = RetimeWrapper_160_io_out;
  assign RetimeWrapper_161_io_flow = 1'h1;
  assign RetimeWrapper_161_io_in = x3503_done;
  assign RetimeWrapper_161_clock = clock;
  assign RetimeWrapper_161_reset = reset;
  assign _T_8703 = RetimeWrapper_161_io_out;
  assign RetimeWrapper_162_io_flow = 1'h1;
  assign RetimeWrapper_162_io_in = x3503_done;
  assign RetimeWrapper_162_clock = clock;
  assign RetimeWrapper_162_reset = reset;
  assign _T_8709 = RetimeWrapper_162_io_out;
  assign RetimeWrapper_163_io_flow = 1'h1;
  assign RetimeWrapper_163_io_in = x3514_done;
  assign RetimeWrapper_163_clock = clock;
  assign RetimeWrapper_163_reset = reset;
  assign _T_8715 = RetimeWrapper_163_io_out;
  assign RetimeWrapper_164_io_flow = 1'h1;
  assign RetimeWrapper_164_io_in = x3503_done;
  assign RetimeWrapper_164_clock = clock;
  assign RetimeWrapper_164_reset = reset;
  assign _T_8721 = RetimeWrapper_164_io_out;
  assign RetimeWrapper_165_io_flow = 1'h1;
  assign RetimeWrapper_165_io_in = x3514_done;
  assign RetimeWrapper_165_clock = clock;
  assign RetimeWrapper_165_reset = reset;
  assign _T_8727 = RetimeWrapper_165_io_out;
  assign RetimeWrapper_166_io_flow = 1'h1;
  assign RetimeWrapper_166_io_in = x3301_done;
  assign RetimeWrapper_166_clock = clock;
  assign RetimeWrapper_166_reset = reset;
  assign _T_8733 = RetimeWrapper_166_io_out;
  assign RetimeWrapper_167_io_flow = 1'h1;
  assign RetimeWrapper_167_io_in = x3428_done;
  assign RetimeWrapper_167_clock = clock;
  assign RetimeWrapper_167_reset = reset;
  assign _T_8739 = RetimeWrapper_167_io_out;
  assign RetimeWrapper_168_io_flow = 1'h1;
  assign RetimeWrapper_168_io_in = x3503_done;
  assign RetimeWrapper_168_clock = clock;
  assign RetimeWrapper_168_reset = reset;
  assign _T_8745 = RetimeWrapper_168_io_out;
  assign RetimeWrapper_169_io_flow = 1'h1;
  assign RetimeWrapper_169_io_in = x3301_done;
  assign RetimeWrapper_169_clock = clock;
  assign RetimeWrapper_169_reset = reset;
  assign _T_8751 = RetimeWrapper_169_io_out;
  assign RetimeWrapper_170_io_flow = 1'h1;
  assign RetimeWrapper_170_io_in = x3428_done;
  assign RetimeWrapper_170_clock = clock;
  assign RetimeWrapper_170_reset = reset;
  assign _T_8757 = RetimeWrapper_170_io_out;
  assign RetimeWrapper_171_io_flow = 1'h1;
  assign RetimeWrapper_171_io_in = x3503_done;
  assign RetimeWrapper_171_clock = clock;
  assign RetimeWrapper_171_reset = reset;
  assign _T_8763 = RetimeWrapper_171_io_out;
  assign RetimeWrapper_172_io_flow = 1'h1;
  assign RetimeWrapper_172_io_in = x3428_done;
  assign RetimeWrapper_172_clock = clock;
  assign RetimeWrapper_172_reset = reset;
  assign _T_8769 = RetimeWrapper_172_io_out;
  assign RetimeWrapper_173_io_flow = 1'h1;
  assign RetimeWrapper_173_io_in = x3503_done;
  assign RetimeWrapper_173_clock = clock;
  assign RetimeWrapper_173_reset = reset;
  assign _T_8775 = RetimeWrapper_173_io_out;
  assign RetimeWrapper_174_io_flow = 1'h1;
  assign RetimeWrapper_174_io_in = x3428_done;
  assign RetimeWrapper_174_clock = clock;
  assign RetimeWrapper_174_reset = reset;
  assign _T_8781 = RetimeWrapper_174_io_out;
  assign RetimeWrapper_175_io_flow = 1'h1;
  assign RetimeWrapper_175_io_in = x3503_done;
  assign RetimeWrapper_175_clock = clock;
  assign RetimeWrapper_175_reset = reset;
  assign _T_8787 = RetimeWrapper_175_io_out;
  assign _T_8821_0_addr_0 = x3474_rVec_0_addr_0;
  assign _T_8821_0_en = x3474_rVec_0_en;
  assign _T_8821_1_addr_0 = x3474_rVec_1_addr_0;
  assign _T_8821_1_en = x3474_rVec_1_en;
  assign _T_8821_2_addr_0 = x3474_rVec_2_addr_0;
  assign _T_8821_2_en = x3474_rVec_2_en;
  assign _T_8821_3_addr_0 = x3474_rVec_3_addr_0;
  assign _T_8821_3_en = x3474_rVec_3_en;
  assign x3474_0_number = x3159_0_io_output_data_8;
  assign x3474_1_number = x3159_0_io_output_data_9;
  assign x3474_2_number = x3159_0_io_output_data_10;
  assign x3474_3_number = x3159_0_io_output_data_11;
  assign _T_8871_0_addr_0 = x3479_rVec_0_addr_0;
  assign _T_8871_0_en = x3479_rVec_0_en;
  assign _T_8871_1_addr_0 = x3479_rVec_1_addr_0;
  assign _T_8871_1_en = x3479_rVec_1_en;
  assign _T_8871_2_addr_0 = x3479_rVec_2_addr_0;
  assign _T_8871_2_en = x3479_rVec_2_en;
  assign _T_8871_3_addr_0 = x3479_rVec_3_addr_0;
  assign _T_8871_3_en = x3479_rVec_3_en;
  assign x3479_0_number = x3161_0_io_output_data_4;
  assign x3479_1_number = x3161_0_io_output_data_5;
  assign x3479_2_number = x3161_0_io_output_data_6;
  assign x3479_3_number = x3161_0_io_output_data_7;
  assign _T_8899_number = _T_8913[31:0];
  assign _T_8915_number = _T_8933;
  assign _T_8926 = _T_8931;
  assign _T_8928 = _T_8926;
  assign _T_8930 = _T_8932;
  assign _T_8935_number = _T_8949[31:0];
  assign _T_8951_number = _T_8969;
  assign _T_8962 = _T_8967;
  assign _T_8964 = _T_8962;
  assign _T_8966 = _T_8968;
  assign _T_8971_number = _T_8985[31:0];
  assign _T_8987_number = _T_9005;
  assign _T_8998 = _T_9003;
  assign _T_9000 = _T_8998;
  assign _T_9002 = _T_9004;
  assign _T_9007_number = _T_9021[31:0];
  assign _T_9023_number = _T_9041;
  assign _T_9034 = _T_9039;
  assign _T_9036 = _T_9034;
  assign _T_9038 = _T_9040;
  assign _T_9043_number = _T_9075;
  assign _T_9045_number = _T_9060;
  assign _T_9047_number = _T_9073;
  assign _T_9051 = _T_9056;
  assign _T_9053 = _T_9051;
  assign _T_9055 = _T_9059;
  assign _T_9064 = _T_9069;
  assign _T_9066 = _T_9064;
  assign _T_9068 = _T_9072;
  assign _T_9077_number = _T_9095;
  assign _T_9087 = _T_9092;
  assign _T_9089 = _T_9087;
  assign _T_9091 = _T_9094;
  assign _T_9099_number = _T_9131;
  assign _T_9101_number = _T_9116;
  assign _T_9103_number = _T_9129;
  assign _T_9107 = _T_9112;
  assign _T_9109 = _T_9107;
  assign _T_9111 = _T_9115;
  assign _T_9120 = _T_9125;
  assign _T_9122 = _T_9120;
  assign _T_9124 = _T_9128;
  assign _T_9133_number = _T_9151;
  assign _T_9143 = _T_9148;
  assign _T_9145 = _T_9143;
  assign _T_9147 = _T_9150;
  assign _T_9155_number = _T_9187;
  assign _T_9157_number = _T_9172;
  assign _T_9159_number = _T_9185;
  assign _T_9163 = _T_9168;
  assign _T_9165 = _T_9163;
  assign _T_9167 = _T_9171;
  assign _T_9176 = _T_9181;
  assign _T_9178 = _T_9176;
  assign _T_9180 = _T_9184;
  assign _T_9189_number = _T_9207;
  assign _T_9199 = _T_9204;
  assign _T_9201 = _T_9199;
  assign _T_9203 = _T_9206;
  assign _T_9217_number = _T_9227;
  assign _T_9227 = b1520_number;
  assign _T_9244_number = _T_9276;
  assign _T_9246_number = _T_9261;
  assign _T_9252 = _T_9257;
  assign _T_9254 = _T_9252;
  assign _T_9256 = _T_9260;
  assign _T_9278_number = _T_9296;
  assign _T_9288 = _T_9293;
  assign _T_9290 = _T_9288;
  assign _T_9292 = _T_9295;
  assign RetimeWrapper_176_io_flow = 1'h1;
  assign RetimeWrapper_176_io_in = x3430_wren;
  assign RetimeWrapper_176_clock = clock;
  assign RetimeWrapper_176_reset = reset;
  assign _T_9309 = RetimeWrapper_176_io_out;
  assign RetimeWrapper_177_io_flow = 1'h1;
  assign RetimeWrapper_177_io_in = reset;
  assign RetimeWrapper_177_clock = clock;
  assign RetimeWrapper_177_reset = reset;
  assign _T_9316 = RetimeWrapper_177_io_out;
  assign RetimeWrapper_178_io_flow = _T_9320;
  assign RetimeWrapper_178_io_in = _T_9336;
  assign RetimeWrapper_178_clock = clock;
  assign RetimeWrapper_178_reset = reset;
  assign _T_9341 = RetimeWrapper_178_io_out;
  assign RetimeWrapper_179_io_flow = _T_9320;
  assign RetimeWrapper_179_io_in = x3364_ctr_trivial;
  assign RetimeWrapper_179_clock = clock;
  assign RetimeWrapper_179_reset = reset;
  assign _T_9350 = RetimeWrapper_179_io_out;
  assign RetimeWrapper_180_io_flow = 1'h1;
  assign RetimeWrapper_180_io_in = x3364_ctr_trivial;
  assign RetimeWrapper_180_clock = clock;
  assign RetimeWrapper_180_reset = reset;
  assign _T_9382 = RetimeWrapper_180_io_out;
  assign RetimeWrapper_181_io_flow = 1'h1;
  assign RetimeWrapper_181_io_in = x3363_sm_io_output_stageEnable_0;
  assign RetimeWrapper_181_clock = clock;
  assign RetimeWrapper_181_reset = reset;
  assign _T_9390 = RetimeWrapper_181_io_out;
  assign RetimeWrapper_182_io_flow = 1'h1;
  assign RetimeWrapper_182_io_in = _T_9393;
  assign RetimeWrapper_182_clock = clock;
  assign RetimeWrapper_182_reset = reset;
  assign _T_9397 = RetimeWrapper_182_io_out;
  assign RetimeWrapper_183_io_flow = 1'h1;
  assign RetimeWrapper_183_io_in = _T_9401;
  assign RetimeWrapper_183_clock = clock;
  assign RetimeWrapper_183_reset = reset;
  assign _T_9405 = RetimeWrapper_183_io_out;
  assign RetimeWrapper_184_io_flow = 1'h1;
  assign RetimeWrapper_184_io_in = x3363_sm_io_output_rst_en;
  assign RetimeWrapper_184_clock = clock;
  assign RetimeWrapper_184_reset = reset;
  assign _T_9414 = RetimeWrapper_184_io_out;
  assign RetimeWrapper_185_io_flow = 1'h1;
  assign RetimeWrapper_185_io_in = x3363_sm_io_output_stageEnable_1;
  assign RetimeWrapper_185_clock = clock;
  assign RetimeWrapper_185_reset = reset;
  assign _T_9420 = RetimeWrapper_185_io_out;
  assign RetimeWrapper_186_io_flow = 1'h1;
  assign RetimeWrapper_186_io_in = _T_9423;
  assign RetimeWrapper_186_clock = clock;
  assign RetimeWrapper_186_reset = reset;
  assign _T_9427 = RetimeWrapper_186_io_out;
  assign RetimeWrapper_187_io_flow = 1'h1;
  assign RetimeWrapper_187_io_in = x3363_sm_io_output_rst_en;
  assign RetimeWrapper_187_clock = clock;
  assign RetimeWrapper_187_reset = reset;
  assign RetimeWrapper_188_io_flow = 1'h1;
  assign RetimeWrapper_188_io_in = _T_9455;
  assign RetimeWrapper_188_clock = clock;
  assign RetimeWrapper_188_reset = reset;
  assign _T_9459 = RetimeWrapper_188_io_out;
  assign RetimeWrapper_189_io_flow = 1'h1;
  assign RetimeWrapper_189_io_in = x3363_ctr_trivial;
  assign RetimeWrapper_189_clock = clock;
  assign RetimeWrapper_189_reset = reset;
  assign _T_9467 = RetimeWrapper_189_io_out;
  assign RetimeWrapper_190_io_flow = 1'h1;
  assign RetimeWrapper_190_io_in = x3362_done;
  assign RetimeWrapper_190_clock = clock;
  assign RetimeWrapper_190_reset = reset;
  assign _T_9753 = RetimeWrapper_190_io_out;
  assign RetimeWrapper_191_io_flow = 1'h1;
  assign RetimeWrapper_191_io_in = x3350_done;
  assign RetimeWrapper_191_clock = clock;
  assign RetimeWrapper_191_reset = reset;
  assign _T_9759 = RetimeWrapper_191_io_out;
  assign _T_9838_number = _T_9848;
  assign _T_9840_number = _T_9859;
  assign _T_9848 = b1393_number;
  assign _T_9859 = x3348_number;
  assign RetimeWrapper_192_io_flow = 1'h1;
  assign RetimeWrapper_192_io_in = x3363_ctr_trivial;
  assign RetimeWrapper_192_clock = clock;
  assign RetimeWrapper_192_reset = reset;
  assign _T_9899 = RetimeWrapper_192_io_out;
  assign _T_9903_number = _T_9913;
  assign _T_9913 = x3348_number;
  assign _T_9932_number = _T_9942;
  assign _T_9934_number = _T_9953;
  assign _T_9942 = x3351_number;
  assign _T_9953 = b1393_number;
  assign _T_9961_number = _T_9971;
  assign _T_9963_number = _T_9982;
  assign _T_9971 = b1393_number;
  assign _T_9982 = x3353_number;
  assign _T_9991_number = _T_10024;
  assign _T_9993_number = _T_10003;
  assign _T_9995_number = _T_10016;
  assign _T_10003 = _T_10008;
  assign _T_10016 = _T_10021;
  assign _T_10026_number = _T_10040;
  assign _T_10040 = _T_10044;
  assign _T_10086_0_addr_0 = x3438_rVec_0_addr_0;
  assign _T_10086_0_en = x3438_rVec_0_en;
  assign _T_10086_1_addr_0 = x3438_rVec_1_addr_0;
  assign _T_10086_1_en = x3438_rVec_1_en;
  assign _T_10086_2_addr_0 = x3438_rVec_2_addr_0;
  assign _T_10086_2_en = x3438_rVec_2_en;
  assign _T_10086_3_addr_0 = x3438_rVec_3_addr_0;
  assign _T_10086_3_en = x3438_rVec_3_en;
  assign x3438_0_number = x3158_0_io_output_data_8;
  assign x3438_1_number = x3158_0_io_output_data_9;
  assign x3438_2_number = x3158_0_io_output_data_10;
  assign x3438_3_number = x3158_0_io_output_data_11;
  assign _T_10136_0_addr_0 = x3443_rVec_0_addr_0;
  assign _T_10136_0_en = x3443_rVec_0_en;
  assign _T_10136_1_addr_0 = x3443_rVec_1_addr_0;
  assign _T_10136_1_en = x3443_rVec_1_en;
  assign _T_10136_2_addr_0 = x3443_rVec_2_addr_0;
  assign _T_10136_2_en = x3443_rVec_2_en;
  assign _T_10136_3_addr_0 = x3443_rVec_3_addr_0;
  assign _T_10136_3_en = x3443_rVec_3_en;
  assign x3443_0_number = x3160_0_io_output_data_4;
  assign x3443_1_number = x3160_0_io_output_data_5;
  assign x3443_2_number = x3160_0_io_output_data_6;
  assign x3443_3_number = x3160_0_io_output_data_7;
  assign _T_10164_number = _T_10178[31:0];
  assign _T_10180_number = _T_10198;
  assign _T_10191 = _T_10196;
  assign _T_10193 = _T_10191;
  assign _T_10195 = _T_10197;
  assign _T_10200_number = _T_10214[31:0];
  assign _T_10216_number = _T_10234;
  assign _T_10227 = _T_10232;
  assign _T_10229 = _T_10227;
  assign _T_10231 = _T_10233;
  assign _T_10236_number = _T_10250[31:0];
  assign _T_10252_number = _T_10270;
  assign _T_10263 = _T_10268;
  assign _T_10265 = _T_10263;
  assign _T_10267 = _T_10269;
  assign _T_10272_number = _T_10286[31:0];
  assign _T_10288_number = _T_10306;
  assign _T_10299 = _T_10304;
  assign _T_10301 = _T_10299;
  assign _T_10303 = _T_10305;
  assign _T_10308_number = _T_10340;
  assign _T_10310_number = _T_10325;
  assign _T_10312_number = _T_10338;
  assign _T_10316 = _T_10321;
  assign _T_10318 = _T_10316;
  assign _T_10320 = _T_10324;
  assign _T_10329 = _T_10334;
  assign _T_10331 = _T_10329;
  assign _T_10333 = _T_10337;
  assign _T_10342_number = _T_10360;
  assign _T_10352 = _T_10357;
  assign _T_10354 = _T_10352;
  assign _T_10356 = _T_10359;
  assign _T_10364_number = _T_10396;
  assign _T_10366_number = _T_10381;
  assign _T_10368_number = _T_10394;
  assign _T_10372 = _T_10377;
  assign _T_10374 = _T_10372;
  assign _T_10376 = _T_10380;
  assign _T_10385 = _T_10390;
  assign _T_10387 = _T_10385;
  assign _T_10389 = _T_10393;
  assign _T_10398_number = _T_10416;
  assign _T_10408 = _T_10413;
  assign _T_10410 = _T_10408;
  assign _T_10412 = _T_10415;
  assign _T_10420_number = _T_10452;
  assign _T_10422_number = _T_10437;
  assign _T_10424_number = _T_10450;
  assign _T_10428 = _T_10433;
  assign _T_10430 = _T_10428;
  assign _T_10432 = _T_10436;
  assign _T_10441 = _T_10446;
  assign _T_10443 = _T_10441;
  assign _T_10445 = _T_10449;
  assign _T_10454_number = _T_10472;
  assign _T_10464 = _T_10469;
  assign _T_10466 = _T_10464;
  assign _T_10468 = _T_10471;
  assign _T_10482_number = _T_10492;
  assign _T_10492 = b1479_number;
  assign _T_10509_number = _T_10541;
  assign _T_10511_number = _T_10526;
  assign _T_10517 = _T_10522;
  assign _T_10519 = _T_10517;
  assign _T_10521 = _T_10525;
  assign _T_10543_number = _T_10561;
  assign _T_10553 = _T_10558;
  assign _T_10555 = _T_10553;
  assign _T_10557 = _T_10560;
  assign RetimeWrapper_193_io_flow = 1'h1;
  assign RetimeWrapper_193_io_in = x3429_wren;
  assign RetimeWrapper_193_clock = clock;
  assign RetimeWrapper_193_reset = reset;
  assign _T_10574 = RetimeWrapper_193_io_out;
  assign RetimeWrapper_194_io_flow = 1'h1;
  assign RetimeWrapper_194_io_in = reset;
  assign RetimeWrapper_194_clock = clock;
  assign RetimeWrapper_194_reset = reset;
  assign _T_10581 = RetimeWrapper_194_io_out;
  assign _T_10584_number = _T_10594;
  assign _T_10586_number = b1202_chain_read_2;
  assign _T_10594 = _T_10586_number;
  assign _T_10599_number = _T_10600[31:0];
  assign _T_10602_number = _T_10603[31:0];
  assign _T_10605_number = _T_10638;
  assign _T_10607_number = _T_10617;
  assign _T_10609_number = _T_10630;
  assign _T_10617 = _T_10622;
  assign _T_10630 = _T_10635;
  assign _T_10640_number = _T_10654;
  assign _T_10654 = _T_10658;
  assign _T_10660_number = _T_10692;
  assign _T_10662_number = _T_10672;
  assign _T_10664_number = _T_10685;
  assign _T_10672 = _T_10622;
  assign _T_10685 = _T_10690;
  assign _T_10694_number = _T_10708;
  assign _T_10708 = _T_10712;
  assign _T_10718_number = _T_10728;
  assign _T_10728 = x3316_number;
  assign _T_10749_number = _T_10782;
  assign _T_10753_number = _T_10774;
  assign _T_10774 = _T_10779;
  assign _T_10784_number = _T_10798;
  assign _T_10798 = _T_10802;
  assign _T_10809_number = _T_10816;
  assign _T_10818_number = _T_10825;
  assign _T_10827_number = _T_10859;
  assign _T_10829_number = _T_10839;
  assign _T_10831_number = _T_10852;
  assign _T_10839 = _T_10844;
  assign _T_10852 = _T_10857;
  assign _T_10861_number = _T_10875;
  assign _T_10875 = _T_10879;
  assign _T_10881_number = _T_10913;
  assign _T_10883_number = _T_10893;
  assign _T_10885_number = _T_10906;
  assign _T_10893 = _T_10857;
  assign _T_10906 = _T_10844;
  assign _T_10915_number = _T_10929;
  assign _T_10929 = _T_10933;
  assign _T_10935_number = _T_10967;
  assign _T_10937_number = _T_10947;
  assign _T_10939_number = _T_10960;
  assign _T_10947 = _T_10952;
  assign _T_10960 = _T_10965;
  assign _T_10969_number = _T_10983;
  assign _T_10983 = _T_10987;
  assign _T_10989_number = _T_11021;
  assign _T_10991_number = _T_11001;
  assign _T_10993_number = _T_11014;
  assign _T_11001 = _T_10690;
  assign _T_11014 = _T_10635;
  assign _T_11023_number = _T_11037;
  assign _T_11037 = _T_11041;
  assign _T_11043_number = _T_11075;
  assign _T_11045_number = _T_11055;
  assign _T_11047_number = _T_11068;
  assign _T_11055 = _T_11060;
  assign _T_11068 = _T_11073;
  assign _T_11077_number = _T_11091;
  assign _T_11091 = _T_11095;
  assign _T_11103 = _T_11112;
  assign _T_11114_number = _T_11124;
  assign _T_11116_number = io_argIns_2;
  assign _T_11124 = _T_11116_number;
  assign _T_11129_number = _T_11161;
  assign _T_11131_number = _T_11141;
  assign _T_11133_number = _T_11154;
  assign _T_11141 = _T_11146;
  assign _T_11154 = _T_11159;
  assign _T_11163_number = _T_11177;
  assign _T_11177 = _T_11181;
  assign _T_11189 = x3329_number;
  assign _T_11214_0 = x3333;
  assign _T_11228_0 = _T_11202;
  assign x3276 = _T_11250_0;
  assign _T_11243_0 = _T_11240;
  assign _T_11250_0 = x3239_io_out_0;
  assign RetimeWrapper_195_io_flow = 1'h1;
  assign RetimeWrapper_195_io_in = reset;
  assign RetimeWrapper_195_clock = clock;
  assign RetimeWrapper_195_reset = reset;
  assign _T_11263 = RetimeWrapper_195_io_out;
  assign RetimeWrapper_196_io_flow = 1'h1;
  assign RetimeWrapper_196_io_in = reset;
  assign RetimeWrapper_196_clock = clock;
  assign RetimeWrapper_196_reset = reset;
  assign _T_11275 = RetimeWrapper_196_io_out;
  assign RetimeWrapper_197_io_flow = 1'h1;
  assign RetimeWrapper_197_io_in = reset;
  assign RetimeWrapper_197_clock = clock;
  assign RetimeWrapper_197_reset = reset;
  assign _T_11287 = RetimeWrapper_197_io_out;
  assign _T_11291_number = _T_11324;
  assign _T_11293_number = _T_11303;
  assign _T_11295_number = _T_11316;
  assign _T_11303 = _T_11308;
  assign _T_11316 = _T_11321;
  assign _T_11326_number = _T_11340;
  assign _T_11340 = _T_11344;
  assign _T_11352_number = _T_11371;
  assign _T_11371 = x3163_number;
  assign RetimeWrapper_198_io_flow = 1'h1;
  assign RetimeWrapper_198_io_in = reset;
  assign RetimeWrapper_198_clock = clock;
  assign RetimeWrapper_198_reset = reset;
  assign _T_11445 = RetimeWrapper_198_io_out;
  assign RetimeWrapper_199_io_flow = 1'h1;
  assign RetimeWrapper_199_io_in = _T_11466;
  assign RetimeWrapper_199_clock = clock;
  assign RetimeWrapper_199_reset = reset;
  assign _T_11470 = RetimeWrapper_199_io_out;
  assign RetimeWrapper_200_io_flow = 1'h1;
  assign RetimeWrapper_200_io_in = x3426_ctr_trivial;
  assign RetimeWrapper_200_clock = clock;
  assign RetimeWrapper_200_reset = reset;
  assign _T_11478 = RetimeWrapper_200_io_out;
  assign RetimeWrapper_201_io_flow = 1'h1;
  assign RetimeWrapper_201_io_in = x3425_done;
  assign RetimeWrapper_201_clock = clock;
  assign RetimeWrapper_201_reset = reset;
  assign _T_11764 = RetimeWrapper_201_io_out;
  assign RetimeWrapper_202_io_flow = 1'h1;
  assign RetimeWrapper_202_io_in = x3413_done;
  assign RetimeWrapper_202_clock = clock;
  assign RetimeWrapper_202_reset = reset;
  assign _T_11770 = RetimeWrapper_202_io_out;
  assign _T_11849_number = _T_11859;
  assign _T_11851_number = _T_11870;
  assign _T_11859 = b1454_number;
  assign _T_11870 = x3411_number;
  assign RetimeWrapper_203_io_flow = 1'h1;
  assign RetimeWrapper_203_io_in = x3426_ctr_trivial;
  assign RetimeWrapper_203_clock = clock;
  assign RetimeWrapper_203_reset = reset;
  assign _T_11910 = RetimeWrapper_203_io_out;
  assign _T_11914_number = _T_11924;
  assign _T_11924 = x3411_number;
  assign _T_11943_number = _T_11953;
  assign _T_11945_number = _T_11964;
  assign _T_11953 = x3414_number;
  assign _T_11964 = b1454_number;
  assign _T_11972_number = _T_11982;
  assign _T_11974_number = _T_11993;
  assign _T_11982 = b1454_number;
  assign _T_11993 = x3416_number;
  assign _T_12002_number = _T_12035;
  assign _T_12004_number = _T_12014;
  assign _T_12006_number = _T_12027;
  assign _T_12014 = _T_12019;
  assign _T_12027 = _T_12032;
  assign _T_12037_number = _T_12051;
  assign _T_12051 = _T_12055;
  assign x3213 = _T_12084_0;
  assign _T_12077_0 = _T_12074;
  assign _T_12084_0 = x3176_io_out_0;
  assign RetimeWrapper_204_io_flow = 1'h1;
  assign RetimeWrapper_204_io_in = reset;
  assign RetimeWrapper_204_clock = clock;
  assign RetimeWrapper_204_reset = reset;
  assign _T_12097 = RetimeWrapper_204_io_out;
  assign RetimeWrapper_205_io_flow = 1'h1;
  assign RetimeWrapper_205_io_in = reset;
  assign RetimeWrapper_205_clock = clock;
  assign RetimeWrapper_205_reset = reset;
  assign _T_12109 = RetimeWrapper_205_io_out;
  assign RetimeWrapper_206_io_flow = 1'h1;
  assign RetimeWrapper_206_io_in = reset;
  assign RetimeWrapper_206_clock = clock;
  assign RetimeWrapper_206_reset = reset;
  assign _T_12121 = RetimeWrapper_206_io_out;
  assign _T_12126_number = _T_12136;
  assign _T_12128_number = _T_12147;
  assign _T_12136 = x3287_number;
  assign _T_12147 = b1331_number;
  assign _T_12155_number = _T_12165;
  assign _T_12157_number = _T_12176;
  assign _T_12165 = b1331_number;
  assign _T_12176 = x3289_number;
  assign _T_12185_number = _T_12218;
  assign _T_12187_number = _T_12197;
  assign _T_12189_number = _T_12210;
  assign _T_12197 = _T_12202;
  assign _T_12210 = _T_12215;
  assign _T_12220_number = _T_12234;
  assign _T_12234 = _T_12238;
  assign _T_12251_number = _T_12261;
  assign _T_12253_number = _T_12272;
  assign _T_12261 = x3224_number;
  assign _T_12272 = b1270_number;
  assign _T_12280_number = _T_12290;
  assign _T_12282_number = _T_12301;
  assign _T_12290 = b1270_number;
  assign _T_12301 = x3226_number;
  assign _T_12310_number = _T_12343;
  assign _T_12312_number = _T_12322;
  assign _T_12314_number = _T_12335;
  assign _T_12322 = _T_12327;
  assign _T_12335 = _T_12340;
  assign _T_12345_number = _T_12359;
  assign _T_12359 = _T_12363;
  assign x3340 = _T_12392_0;
  assign _T_12385_0 = _T_12382;
  assign _T_12392_0 = x3303_io_out_0;
  assign RetimeWrapper_207_io_flow = 1'h1;
  assign RetimeWrapper_207_io_in = reset;
  assign RetimeWrapper_207_clock = clock;
  assign RetimeWrapper_207_reset = reset;
  assign _T_12405 = RetimeWrapper_207_io_out;
  assign RetimeWrapper_208_io_flow = 1'h1;
  assign RetimeWrapper_208_io_in = reset;
  assign RetimeWrapper_208_clock = clock;
  assign RetimeWrapper_208_reset = reset;
  assign _T_12417 = RetimeWrapper_208_io_out;
  assign RetimeWrapper_209_io_flow = 1'h1;
  assign RetimeWrapper_209_io_in = reset;
  assign RetimeWrapper_209_clock = clock;
  assign RetimeWrapper_209_reset = reset;
  assign _T_12429 = RetimeWrapper_209_io_out;
  assign x3403 = _T_12450_0;
  assign _T_12443_0 = _T_12440;
  assign _T_12450_0 = x3366_io_out_0;
  assign RetimeWrapper_210_io_flow = 1'h1;
  assign RetimeWrapper_210_io_in = reset;
  assign RetimeWrapper_210_clock = clock;
  assign RetimeWrapper_210_reset = reset;
  assign _T_12463 = RetimeWrapper_210_io_out;
  assign RetimeWrapper_211_io_flow = 1'h1;
  assign RetimeWrapper_211_io_in = reset;
  assign RetimeWrapper_211_clock = clock;
  assign RetimeWrapper_211_reset = reset;
  assign _T_12475 = RetimeWrapper_211_io_out;
  assign RetimeWrapper_212_io_flow = 1'h1;
  assign RetimeWrapper_212_io_in = reset;
  assign RetimeWrapper_212_clock = clock;
  assign RetimeWrapper_212_reset = reset;
  assign _T_12487 = RetimeWrapper_212_io_out;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_1682 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_1985 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  _T_2433 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  _T_2448 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  _T_2524 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  _T_2594 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  _T_2664 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  _T_2736 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  _T_2806 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  _T_2821 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  _T_2996 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  _T_3115 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  _T_3746 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  _T_4515 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  _T_4634 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  _T_5389 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  _T_6247 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  _T_8324 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  _T_8339 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  _T_8370 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  _T_8385 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  _T_9330 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  _T_9449 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  _T_11460 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_1682 <= 1'h0;
    end else begin
      _T_1682 <= _T_1679;
    end
    if (reset) begin
      _T_1985 <= 1'h0;
    end else begin
      _T_1985 <= _T_1982;
    end
    if (reset) begin
      _T_2433 <= 1'h0;
    end else begin
      _T_2433 <= _T_2430;
    end
    if (reset) begin
      _T_2448 <= 1'h0;
    end else begin
      _T_2448 <= _T_2445;
    end
    if (reset) begin
      _T_2524 <= 1'h0;
    end else begin
      _T_2524 <= _T_2521;
    end
    if (reset) begin
      _T_2594 <= 1'h0;
    end else begin
      _T_2594 <= _T_2591;
    end
    if (reset) begin
      _T_2664 <= 1'h0;
    end else begin
      _T_2664 <= _T_2661;
    end
    if (reset) begin
      _T_2736 <= 1'h0;
    end else begin
      _T_2736 <= _T_2733;
    end
    if (reset) begin
      _T_2806 <= 1'h0;
    end else begin
      _T_2806 <= _T_2803;
    end
    if (reset) begin
      _T_2821 <= 1'h0;
    end else begin
      _T_2821 <= _T_2818;
    end
    if (reset) begin
      _T_2996 <= 1'h0;
    end else begin
      _T_2996 <= _T_2993;
    end
    if (reset) begin
      _T_3115 <= 1'h0;
    end else begin
      _T_3115 <= _T_3112;
    end
    if (reset) begin
      _T_3746 <= 1'h0;
    end else begin
      _T_3746 <= _T_3743;
    end
    if (reset) begin
      _T_4515 <= 1'h0;
    end else begin
      _T_4515 <= _T_4512;
    end
    if (reset) begin
      _T_4634 <= 1'h0;
    end else begin
      _T_4634 <= _T_4631;
    end
    if (reset) begin
      _T_5389 <= 1'h0;
    end else begin
      _T_5389 <= _T_5386;
    end
    if (reset) begin
      _T_6247 <= 1'h0;
    end else begin
      _T_6247 <= _T_6244;
    end
    if (reset) begin
      _T_8324 <= 1'h0;
    end else begin
      _T_8324 <= _T_8321;
    end
    if (reset) begin
      _T_8339 <= 1'h0;
    end else begin
      _T_8339 <= _T_8336;
    end
    if (reset) begin
      _T_8370 <= 1'h0;
    end else begin
      _T_8370 <= _T_8367;
    end
    if (reset) begin
      _T_8385 <= 1'h0;
    end else begin
      _T_8385 <= _T_8382;
    end
    if (reset) begin
      _T_9330 <= 1'h0;
    end else begin
      _T_9330 <= _T_9327;
    end
    if (reset) begin
      _T_9449 <= 1'h0;
    end else begin
      _T_9449 <= _T_9446;
    end
    if (reset) begin
      _T_11460 <= 1'h0;
    end else begin
      _T_11460 <= _T_11457;
    end
  end
endmodule
module FF_115(
  input   clock,
  input   reset,
  input   io_in,
  input   io_init,
  input   io_reset,
  output  io_out,
  input   io_enable
);
  wire  d;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire  RetimeWrapper_io_flow;
  wire  RetimeWrapper_io_in;
  wire  RetimeWrapper_io_out;
  wire  _T_11;
  wire  _GEN_0;
  wire  _GEN_1;
  RetimeWrapper RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _GEN_0 = io_reset ? io_init : _T_11;
  assign _GEN_1 = io_enable ? io_in : _GEN_0;
  assign io_out = _T_11;
  assign d = _GEN_1;
  assign RetimeWrapper_io_flow = 1'h1;
  assign RetimeWrapper_io_in = d;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_11 = RetimeWrapper_io_out;
endmodule
module MuxN(
  input  [63:0] io_ins_0_0_addr,
  input         io_ins_0_0_isWr,
  input  [15:0] io_ins_0_0_size,
  input  [63:0] io_ins_1_0_addr,
  input         io_ins_1_0_isWr,
  input  [15:0] io_ins_1_0_size,
  input         io_sel,
  output [63:0] io_out_0_addr,
  output        io_out_0_isWr,
  output [15:0] io_out_0_size
);
  wire [15:0] _GEN_0_0_size;
  wire [63:0] _GEN_4;
  wire  _GEN_5;
  wire [15:0] _GEN_7;
  wire  _GEN_2_0_isWr;
  wire [63:0] _GEN_3_0_addr;
  assign _GEN_4 = io_sel ? io_ins_1_0_addr : io_ins_0_0_addr;
  assign _GEN_5 = io_sel ? io_ins_1_0_isWr : io_ins_0_0_isWr;
  assign _GEN_7 = io_sel ? io_ins_1_0_size : io_ins_0_0_size;
  assign io_out_0_addr = _GEN_3_0_addr;
  assign io_out_0_isWr = _GEN_2_0_isWr;
  assign io_out_0_size = _GEN_0_0_size;
  assign _GEN_0_0_size = _GEN_7;
  assign _GEN_2_0_isWr = _GEN_5;
  assign _GEN_3_0_addr = _GEN_4;
endmodule
module MuxNPipe(
  input  [63:0] io_ins_0_0_addr,
  input         io_ins_0_0_isWr,
  input  [15:0] io_ins_0_0_size,
  input  [63:0] io_ins_1_0_addr,
  input         io_ins_1_0_isWr,
  input  [15:0] io_ins_1_0_size,
  input         io_sel,
  output [63:0] io_out_0_addr,
  output        io_out_0_isWr,
  output [15:0] io_out_0_size
);
  wire [63:0] _T_103_0_0_addr;
  wire  _T_103_0_0_isWr;
  wire [15:0] _T_103_0_0_size;
  wire [63:0] _T_103_1_0_addr;
  wire  _T_103_1_0_isWr;
  wire [15:0] _T_103_1_0_size;
  wire [63:0] MuxN_io_ins_0_0_addr;
  wire  MuxN_io_ins_0_0_isWr;
  wire [15:0] MuxN_io_ins_0_0_size;
  wire [63:0] MuxN_io_ins_1_0_addr;
  wire  MuxN_io_ins_1_0_isWr;
  wire [15:0] MuxN_io_ins_1_0_size;
  wire  MuxN_io_sel;
  wire [63:0] MuxN_io_out_0_addr;
  wire  MuxN_io_out_0_isWr;
  wire [15:0] MuxN_io_out_0_size;
  MuxN MuxN (
    .io_ins_0_0_addr(MuxN_io_ins_0_0_addr),
    .io_ins_0_0_isWr(MuxN_io_ins_0_0_isWr),
    .io_ins_0_0_size(MuxN_io_ins_0_0_size),
    .io_ins_1_0_addr(MuxN_io_ins_1_0_addr),
    .io_ins_1_0_isWr(MuxN_io_ins_1_0_isWr),
    .io_ins_1_0_size(MuxN_io_ins_1_0_size),
    .io_sel(MuxN_io_sel),
    .io_out_0_addr(MuxN_io_out_0_addr),
    .io_out_0_isWr(MuxN_io_out_0_isWr),
    .io_out_0_size(MuxN_io_out_0_size)
  );
  assign io_out_0_addr = MuxN_io_out_0_addr;
  assign io_out_0_isWr = MuxN_io_out_0_isWr;
  assign io_out_0_size = MuxN_io_out_0_size;
  assign _T_103_0_0_addr = io_ins_0_0_addr;
  assign _T_103_0_0_isWr = io_ins_0_0_isWr;
  assign _T_103_0_0_size = io_ins_0_0_size;
  assign _T_103_1_0_addr = io_ins_1_0_addr;
  assign _T_103_1_0_isWr = io_ins_1_0_isWr;
  assign _T_103_1_0_size = io_ins_1_0_size;
  assign MuxN_io_ins_0_0_addr = _T_103_0_0_addr;
  assign MuxN_io_ins_0_0_isWr = _T_103_0_0_isWr;
  assign MuxN_io_ins_0_0_size = _T_103_0_0_size;
  assign MuxN_io_ins_1_0_addr = _T_103_1_0_addr;
  assign MuxN_io_ins_1_0_isWr = _T_103_1_0_isWr;
  assign MuxN_io_ins_1_0_size = _T_103_1_0_size;
  assign MuxN_io_sel = io_sel;
endmodule
module FIFOArbiter(
  input         clock,
  input         reset,
  output [63:0] io_fifo_0_enq_0_addr,
  output        io_fifo_0_enq_0_isWr,
  output [15:0] io_fifo_0_enq_0_size,
  output        io_fifo_0_enqVld,
  input  [63:0] io_fifo_0_deq_0_addr,
  input         io_fifo_0_deq_0_isWr,
  input  [15:0] io_fifo_0_deq_0_size,
  output        io_fifo_0_deqVld,
  input         io_fifo_0_full,
  input         io_fifo_0_empty,
  input         io_fifo_0_almostEmpty,
  input  [63:0] io_fifo_1_deq_0_addr,
  input         io_fifo_1_deq_0_isWr,
  input  [15:0] io_fifo_1_deq_0_size,
  output        io_fifo_1_deqVld,
  input         io_fifo_1_empty,
  input  [63:0] io_enq_0_0_addr,
  input         io_enq_0_0_isWr,
  input  [15:0] io_enq_0_0_size,
  input         io_enqVld_0,
  output        io_full_0,
  output [63:0] io_deq_0_addr,
  output        io_deq_0_isWr,
  output [15:0] io_deq_0_size,
  input         io_deqVld,
  output        io_deqReady,
  output        io_empty,
  output        io_tag
);
  wire  tagFF_clock;
  wire  tagFF_reset;
  wire  tagFF_io_in;
  wire  tagFF_io_init;
  wire  tagFF_io_reset;
  wire  tagFF_io_out;
  wire  tagFF_io_enable;
  wire  tag;
  wire  _T_173;
  wire  _T_174;
  wire  _T_179;
  wire  _T_181;
  wire  _T_182;
  wire  _T_183;
  wire  _T_184;
  wire  _T_185;
  wire  _T_188;
  wire  _T_190;
  wire  _T_191;
  wire  _T_192;
  wire  _T_193;
  wire  _T_206_0;
  wire  _T_211_0;
  wire  _T_221;
  wire  _T_226;
  wire  _T_227;
  wire  _T_228;
  wire [63:0] MuxNPipe_io_ins_0_0_addr;
  wire  MuxNPipe_io_ins_0_0_isWr;
  wire [15:0] MuxNPipe_io_ins_0_0_size;
  wire [63:0] MuxNPipe_io_ins_1_0_addr;
  wire  MuxNPipe_io_ins_1_0_isWr;
  wire [15:0] MuxNPipe_io_ins_1_0_size;
  wire  MuxNPipe_io_sel;
  wire [63:0] MuxNPipe_io_out_0_addr;
  wire  MuxNPipe_io_out_0_isWr;
  wire [15:0] MuxNPipe_io_out_0_size;
  wire [63:0] _T_247_0_0_addr;
  wire  _T_247_0_0_isWr;
  wire [15:0] _T_247_0_0_size;
  wire [63:0] _T_247_1_0_addr;
  wire  _T_247_1_0_isWr;
  wire [15:0] _T_247_1_0_size;
  wire  _T_288;
  FF_115 tagFF (
    .clock(tagFF_clock),
    .reset(tagFF_reset),
    .io_in(tagFF_io_in),
    .io_init(tagFF_io_init),
    .io_reset(tagFF_io_reset),
    .io_out(tagFF_io_out),
    .io_enable(tagFF_io_enable)
  );
  MuxNPipe MuxNPipe (
    .io_ins_0_0_addr(MuxNPipe_io_ins_0_0_addr),
    .io_ins_0_0_isWr(MuxNPipe_io_ins_0_0_isWr),
    .io_ins_0_0_size(MuxNPipe_io_ins_0_0_size),
    .io_ins_1_0_addr(MuxNPipe_io_ins_1_0_addr),
    .io_ins_1_0_isWr(MuxNPipe_io_ins_1_0_isWr),
    .io_ins_1_0_size(MuxNPipe_io_ins_1_0_size),
    .io_sel(MuxNPipe_io_sel),
    .io_out_0_addr(MuxNPipe_io_out_0_addr),
    .io_out_0_isWr(MuxNPipe_io_out_0_isWr),
    .io_out_0_size(MuxNPipe_io_out_0_size)
  );
  assign tag = tagFF_io_out;
  assign _T_173 = tag == 1'h0;
  assign _T_174 = io_deqVld & _T_173;
  assign _T_179 = io_deqVld & tag;
  assign _T_181 = io_fifo_0_empty & io_fifo_1_empty;
  assign _T_182 = _T_181 & io_enqVld_0;
  assign _T_183 = io_deqVld | _T_182;
  assign _T_184 = ~ io_enqVld_0;
  assign _T_185 = _T_184 & io_fifo_0_empty;
  assign _T_188 = _T_173 & io_deqVld;
  assign _T_190 = _T_188 & _T_184;
  assign _T_191 = _T_190 & io_fifo_0_almostEmpty;
  assign _T_192 = _T_185 | _T_191;
  assign _T_193 = ~ _T_192;
  assign _T_211_0 = _T_181 ? io_enqVld_0 : _T_206_0;
  assign _T_221 = _T_211_0 ? 1'h0 : 1'h1;
  assign _T_226 = tag ? io_fifo_1_empty : 1'h0;
  assign _T_227 = 1'h0 == tag;
  assign _T_228 = _T_227 ? io_fifo_0_empty : _T_226;
  assign _T_288 = ~ _T_228;
  assign io_fifo_0_enq_0_addr = io_enq_0_0_addr;
  assign io_fifo_0_enq_0_isWr = io_enq_0_0_isWr;
  assign io_fifo_0_enq_0_size = io_enq_0_0_size;
  assign io_fifo_0_enqVld = io_enqVld_0;
  assign io_fifo_0_deqVld = _T_174;
  assign io_fifo_1_deqVld = _T_179;
  assign io_full_0 = io_fifo_0_full;
  assign io_deq_0_addr = MuxNPipe_io_out_0_addr;
  assign io_deq_0_isWr = MuxNPipe_io_out_0_isWr;
  assign io_deq_0_size = MuxNPipe_io_out_0_size;
  assign io_deqReady = _T_288;
  assign io_empty = _T_228;
  assign io_tag = tag;
  assign tagFF_io_in = _T_221;
  assign tagFF_io_init = 1'h0;
  assign tagFF_io_reset = 1'h0;
  assign tagFF_io_enable = _T_183;
  assign tagFF_clock = clock;
  assign tagFF_reset = reset;
  assign _T_206_0 = _T_193;
  assign MuxNPipe_io_ins_0_0_addr = _T_247_0_0_addr;
  assign MuxNPipe_io_ins_0_0_isWr = _T_247_0_0_isWr;
  assign MuxNPipe_io_ins_0_0_size = _T_247_0_0_size;
  assign MuxNPipe_io_ins_1_0_addr = _T_247_1_0_addr;
  assign MuxNPipe_io_ins_1_0_isWr = _T_247_1_0_isWr;
  assign MuxNPipe_io_ins_1_0_size = _T_247_1_0_size;
  assign MuxNPipe_io_sel = tag;
  assign _T_247_0_0_addr = io_fifo_0_deq_0_addr;
  assign _T_247_0_0_isWr = io_fifo_0_deq_0_isWr;
  assign _T_247_0_0_size = io_fifo_0_deq_0_size;
  assign _T_247_1_0_addr = io_fifo_1_deq_0_addr;
  assign _T_247_1_0_isWr = io_fifo_1_deq_0_isWr;
  assign _T_247_1_0_size = io_fifo_1_deq_0_size;
endmodule
module RetimeWrapper_561(
  input        clock,
  input        reset,
  input  [8:0] io_in,
  output [8:0] io_out
);
  wire [8:0] sr_out;
  wire [8:0] sr_in;
  wire  sr_flow;
  wire  sr_reset;
  wire  sr_clock;
  RetimeShiftRegister #(.WIDTH(9), .STAGES(1)) sr (
    .out(sr_out),
    .in(sr_in),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out;
  assign sr_in = io_in;
  assign sr_flow = 1'h1;
  assign sr_reset = reset;
  assign sr_clock = clock;
endmodule
module FF_116(
  input        clock,
  input        reset,
  input  [8:0] io_in,
  output [8:0] io_out,
  input        io_enable
);
  wire [8:0] d;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire [8:0] RetimeWrapper_io_in;
  wire [8:0] RetimeWrapper_io_out;
  wire [8:0] _T_11;
  wire [8:0] _GEN_1;
  RetimeWrapper_561 RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _GEN_1 = io_enable ? io_in : _T_11;
  assign io_out = _T_11;
  assign d = _GEN_1;
  assign RetimeWrapper_io_in = d;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_11 = RetimeWrapper_io_out;
endmodule
module UpDownCtr(
  input        clock,
  input        reset,
  input  [8:0] io_strideInc,
  input  [8:0] io_strideDec,
  input        io_inc,
  input        io_dec,
  output [8:0] io_out,
  output [8:0] io_nextInc,
  output [8:0] io_nextDec
);
  wire  reg$_clock;
  wire  reg$_reset;
  wire [8:0] reg$_io_in;
  wire [8:0] reg$_io_out;
  wire  reg$_io_enable;
  wire  _T_16;
  wire [8:0] incval;
  wire [8:0] decval;
  wire [9:0] _T_20;
  wire [9:0] _T_21;
  wire [8:0] incr;
  wire [9:0] _T_22;
  wire [8:0] newval;
  wire [9:0] _T_27;
  wire [8:0] _T_28;
  wire [9:0] _T_29;
  wire [9:0] _T_30;
  wire [8:0] _T_31;
  FF_116 reg$ (
    .clock(reg$_clock),
    .reset(reg$_reset),
    .io_in(reg$_io_in),
    .io_out(reg$_io_out),
    .io_enable(reg$_io_enable)
  );
  assign _T_16 = io_inc | io_dec;
  assign incval = io_inc ? io_strideInc : 9'h0;
  assign decval = io_dec ? io_strideDec : 9'h0;
  assign _T_20 = incval - decval;
  assign _T_21 = $unsigned(_T_20);
  assign incr = _T_21[8:0];
  assign _T_22 = reg$_io_out + incr;
  assign newval = _T_22[8:0];
  assign _T_27 = reg$_io_out + io_strideInc;
  assign _T_28 = _T_27[8:0];
  assign _T_29 = reg$_io_out - io_strideDec;
  assign _T_30 = $unsigned(_T_29);
  assign _T_31 = _T_30[8:0];
  assign io_out = reg$_io_out;
  assign io_nextInc = _T_28;
  assign io_nextDec = _T_31;
  assign reg$_io_in = newval;
  assign reg$_io_enable = _T_16;
  assign reg$_clock = clock;
  assign reg$_reset = reset;
endmodule
module Counter_7(
  input        clock,
  input        reset,
  input  [8:0] io_max,
  output [8:0] io_out,
  output [8:0] io_next,
  input        io_enable,
  output       io_done
);
  wire  reg$_clock;
  wire  reg$_reset;
  wire [8:0] reg$_io_in;
  wire [8:0] reg$_io_out;
  wire  reg$_io_enable;
  wire [9:0] count;
  wire [10:0] _T_13;
  wire [9:0] newval;
  wire [9:0] _GEN_1;
  wire  isMax;
  wire [9:0] next;
  wire  _T_15;
  FF_116 reg$ (
    .clock(reg$_clock),
    .reset(reg$_reset),
    .io_in(reg$_io_in),
    .io_out(reg$_io_out),
    .io_enable(reg$_io_enable)
  );
  assign count = {1'h0,reg$_io_out};
  assign _T_13 = count + 10'h1;
  assign newval = _T_13[9:0];
  assign _GEN_1 = {{1'd0}, io_max};
  assign isMax = newval >= _GEN_1;
  assign next = isMax ? 10'h0 : newval;
  assign _T_15 = io_enable & isMax;
  assign io_out = count[8:0];
  assign io_next = next[8:0];
  assign io_done = _T_15;
  assign reg$_io_in = next[8:0];
  assign reg$_io_enable = io_enable;
  assign reg$_clock = clock;
  assign reg$_reset = reset;
endmodule
module Depulser(
  input   clock,
  input   reset,
  input   io_in,
  input   io_rst,
  output  io_out
);
  wire  r_clock;
  wire  r_reset;
  wire  r_io_in;
  wire  r_io_init;
  wire  r_io_reset;
  wire  r_io_out;
  wire  r_io_enable;
  wire  _T_6;
  wire  _T_8;
  FF_115 r (
    .clock(r_clock),
    .reset(r_reset),
    .io_in(r_io_in),
    .io_init(r_io_init),
    .io_reset(r_io_reset),
    .io_out(r_io_out),
    .io_enable(r_io_enable)
  );
  assign _T_6 = io_rst ? 1'h0 : io_in;
  assign _T_8 = io_in | io_rst;
  assign io_out = r_io_out;
  assign r_io_in = _T_6;
  assign r_io_init = 1'h0;
  assign r_io_reset = 1'h0;
  assign r_io_enable = _T_8;
  assign r_clock = clock;
  assign r_reset = reset;
endmodule
module CounterCore(
  input        clock,
  input        reset,
  output [8:0] io_out,
  output [8:0] io_next,
  input        io_enable,
  output       io_done,
  input  [8:0] io_config_max
);
  wire  counter_clock;
  wire  counter_reset;
  wire [8:0] counter_io_max;
  wire [8:0] counter_io_out;
  wire [8:0] counter_io_next;
  wire  counter_io_enable;
  wire  counter_io_done;
  wire  depulser_clock;
  wire  depulser_reset;
  wire  depulser_io_in;
  wire  depulser_io_rst;
  wire  depulser_io_out;
  Counter_7 counter (
    .clock(counter_clock),
    .reset(counter_reset),
    .io_max(counter_io_max),
    .io_out(counter_io_out),
    .io_next(counter_io_next),
    .io_enable(counter_io_enable),
    .io_done(counter_io_done)
  );
  Depulser depulser (
    .clock(depulser_clock),
    .reset(depulser_reset),
    .io_in(depulser_io_in),
    .io_rst(depulser_io_rst),
    .io_out(depulser_io_out)
  );
  assign io_out = counter_io_out;
  assign io_next = counter_io_next;
  assign io_done = counter_io_done;
  assign counter_io_max = io_config_max;
  assign counter_io_enable = io_enable;
  assign counter_clock = clock;
  assign counter_reset = reset;
  assign depulser_io_in = counter_io_done;
  assign depulser_io_rst = 1'h0;
  assign depulser_clock = clock;
  assign depulser_reset = reset;
endmodule
module CounterChainCore(
  input        clock,
  input        reset,
  output [8:0] io_out_0,
  output [8:0] io_out_1,
  output [8:0] io_next_1,
  input        io_enable_0,
  input        io_enable_1,
  output       io_done_0,
  input        io_config_chain_0
);
  wire  counters_0_clock;
  wire  counters_0_reset;
  wire [8:0] counters_0_io_out;
  wire [8:0] counters_0_io_next;
  wire  counters_0_io_enable;
  wire  counters_0_io_done;
  wire [8:0] counters_0_io_config_max;
  wire  counters_1_clock;
  wire  counters_1_reset;
  wire [8:0] counters_1_io_out;
  wire [8:0] counters_1_io_next;
  wire  counters_1_io_enable;
  wire  counters_1_io_done;
  wire [8:0] counters_1_io_config_max;
  wire  _T_69;
  CounterCore counters_0 (
    .clock(counters_0_clock),
    .reset(counters_0_reset),
    .io_out(counters_0_io_out),
    .io_next(counters_0_io_next),
    .io_enable(counters_0_io_enable),
    .io_done(counters_0_io_done),
    .io_config_max(counters_0_io_config_max)
  );
  CounterCore counters_1 (
    .clock(counters_1_clock),
    .reset(counters_1_reset),
    .io_out(counters_1_io_out),
    .io_next(counters_1_io_next),
    .io_enable(counters_1_io_enable),
    .io_done(counters_1_io_done),
    .io_config_max(counters_1_io_config_max)
  );
  assign _T_69 = io_config_chain_0 ? counters_0_io_done : io_enable_1;
  assign io_out_0 = counters_0_io_out;
  assign io_out_1 = counters_1_io_out;
  assign io_next_1 = counters_1_io_next;
  assign io_done_0 = counters_0_io_done;
  assign counters_0_io_enable = io_enable_0;
  assign counters_0_io_config_max = 9'h1;
  assign counters_0_clock = clock;
  assign counters_0_reset = reset;
  assign counters_1_io_enable = _T_69;
  assign counters_1_io_config_max = 9'h100;
  assign counters_1_clock = clock;
  assign counters_1_reset = reset;
endmodule
module SRAM_10(
  input         clock,
  input         reset,
  input  [7:0]  io_raddr,
  input         io_wen,
  input  [7:0]  io_waddr,
  input  [63:0] io_wdata_addr,
  input         io_wdata_isWr,
  input  [15:0] io_wdata_size,
  output [63:0] io_rdata_addr,
  output        io_rdata_isWr,
  output [15:0] io_rdata_size
);
  wire [81:0] SRAMVerilogAWS_rdata;
  wire [81:0] SRAMVerilogAWS_wdata;
  wire  SRAMVerilogAWS_flow;
  wire  SRAMVerilogAWS_wen;
  wire  SRAMVerilogAWS_waddrEn;
  wire  SRAMVerilogAWS_raddrEn;
  wire [7:0] SRAMVerilogAWS_waddr;
  wire [7:0] SRAMVerilogAWS_raddr;
  wire  SRAMVerilogAWS_clk;
  wire [16:0] _T_6;
  wire [64:0] _T_7;
  wire [81:0] _T_8;
  wire  _T_11;
  wire  _T_12;
  reg  _T_15;
  reg [31:0] _RAND_0;
  reg [81:0] _T_21;
  reg [95:0] _RAND_1;
  wire [81:0] _T_22;
  wire [63:0] _T_24_addr;
  wire  _T_24_isWr;
  wire [15:0] _T_24_size;
  wire [81:0] _T_26;
  wire [15:0] _T_27;
  wire  _T_29;
  wire [63:0] _T_30;
  SRAMVerilogAWS #(.DWIDTH(82), .WORDS(256), .AWIDTH(8)) SRAMVerilogAWS (
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .flow(SRAMVerilogAWS_flow),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_6 = {1'h0,io_wdata_size};
  assign _T_7 = {io_wdata_addr,io_wdata_isWr};
  assign _T_8 = {_T_7,_T_6};
  assign _T_11 = io_raddr == io_waddr;
  assign _T_12 = io_wen & _T_11;
  assign _T_22 = _T_15 ? _T_21 : SRAMVerilogAWS_rdata;
  assign _T_27 = _T_26[15:0];
  assign _T_29 = _T_26[17];
  assign _T_30 = _T_26[81:18];
  assign io_rdata_addr = _T_24_addr;
  assign io_rdata_isWr = _T_24_isWr;
  assign io_rdata_size = _T_24_size;
  assign SRAMVerilogAWS_wdata = _T_8;
  assign SRAMVerilogAWS_flow = 1'h1;
  assign SRAMVerilogAWS_wen = io_wen;
  assign SRAMVerilogAWS_waddrEn = 1'h1;
  assign SRAMVerilogAWS_raddrEn = 1'h1;
  assign SRAMVerilogAWS_waddr = io_waddr;
  assign SRAMVerilogAWS_raddr = io_raddr;
  assign SRAMVerilogAWS_clk = clock;
  assign _T_24_addr = _T_30;
  assign _T_24_isWr = _T_29;
  assign _T_24_size = _T_27;
  assign _T_26 = _T_22;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_15 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {3{$random}};
  _T_21 = _RAND_1[81:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_15 <= 1'h0;
    end else begin
      _T_15 <= _T_12;
    end
    if (reset) begin
      _T_21 <= 82'h0;
    end else begin
      _T_21 <= _T_8;
    end
  end
endmodule
module MuxN_2(
  input  [63:0] io_ins_0_addr,
  input         io_ins_0_isWr,
  input  [15:0] io_ins_0_size,
  output [63:0] io_out_addr,
  output        io_out_isWr,
  output [15:0] io_out_size
);
  assign io_out_addr = io_ins_0_addr;
  assign io_out_isWr = io_ins_0_isWr;
  assign io_out_size = io_ins_0_size;
endmodule
module FIFOCore(
  input         clock,
  input         reset,
  input  [63:0] io_enq_0_addr,
  input         io_enq_0_isWr,
  input  [15:0] io_enq_0_size,
  input         io_enqVld,
  output [63:0] io_deq_0_addr,
  output        io_deq_0_isWr,
  output [15:0] io_deq_0_size,
  input         io_deqVld,
  output        io_full,
  output        io_empty,
  output        io_almostEmpty
);
  wire  sizeUDC_clock;
  wire  sizeUDC_reset;
  wire [8:0] sizeUDC_io_strideInc;
  wire [8:0] sizeUDC_io_strideDec;
  wire  sizeUDC_io_inc;
  wire  sizeUDC_io_dec;
  wire [8:0] sizeUDC_io_out;
  wire [8:0] sizeUDC_io_nextInc;
  wire [8:0] sizeUDC_io_nextDec;
  wire [9:0] _T_21;
  wire [9:0] _T_22;
  wire [8:0] remainingSlots;
  wire  empty;
  wire  almostEmpty;
  wire  full;
  wire  _T_34;
  wire  writeEn;
  wire  _T_35;
  wire  readEn;
  wire  wptr_clock;
  wire  wptr_reset;
  wire [8:0] wptr_io_out_0;
  wire [8:0] wptr_io_out_1;
  wire [8:0] wptr_io_next_1;
  wire  wptr_io_enable_0;
  wire  wptr_io_enable_1;
  wire  wptr_io_done_0;
  wire  wptr_io_config_chain_0;
  wire  rptr_clock;
  wire  rptr_reset;
  wire [8:0] rptr_io_out_0;
  wire [8:0] rptr_io_out_1;
  wire [8:0] rptr_io_next_1;
  wire  rptr_io_enable_0;
  wire  rptr_io_enable_1;
  wire  rptr_io_done_0;
  wire  rptr_io_config_chain_0;
  wire [8:0] nextHeadLocalAddr;
  wire  mems_0_0_clock;
  wire  mems_0_0_reset;
  wire [7:0] mems_0_0_io_raddr;
  wire  mems_0_0_io_wen;
  wire [7:0] mems_0_0_io_waddr;
  wire [63:0] mems_0_0_io_wdata_addr;
  wire  mems_0_0_io_wdata_isWr;
  wire [15:0] mems_0_0_io_wdata_size;
  wire [63:0] mems_0_0_io_rdata_addr;
  wire  mems_0_0_io_rdata_isWr;
  wire [15:0] mems_0_0_io_rdata_size;
  wire [63:0] wdata_0_addr;
  wire  wdata_0_isWr;
  wire [15:0] wdata_0_size;
  wire [8:0] _T_79;
  wire  _T_81;
  wire  _T_82;
  wire [63:0] MuxN_io_ins_0_addr;
  wire  MuxN_io_ins_0_isWr;
  wire [15:0] MuxN_io_ins_0_size;
  wire [63:0] MuxN_io_out_addr;
  wire  MuxN_io_out_isWr;
  wire [15:0] MuxN_io_out_size;
  UpDownCtr sizeUDC (
    .clock(sizeUDC_clock),
    .reset(sizeUDC_reset),
    .io_strideInc(sizeUDC_io_strideInc),
    .io_strideDec(sizeUDC_io_strideDec),
    .io_inc(sizeUDC_io_inc),
    .io_dec(sizeUDC_io_dec),
    .io_out(sizeUDC_io_out),
    .io_nextInc(sizeUDC_io_nextInc),
    .io_nextDec(sizeUDC_io_nextDec)
  );
  CounterChainCore wptr (
    .clock(wptr_clock),
    .reset(wptr_reset),
    .io_out_0(wptr_io_out_0),
    .io_out_1(wptr_io_out_1),
    .io_next_1(wptr_io_next_1),
    .io_enable_0(wptr_io_enable_0),
    .io_enable_1(wptr_io_enable_1),
    .io_done_0(wptr_io_done_0),
    .io_config_chain_0(wptr_io_config_chain_0)
  );
  CounterChainCore rptr (
    .clock(rptr_clock),
    .reset(rptr_reset),
    .io_out_0(rptr_io_out_0),
    .io_out_1(rptr_io_out_1),
    .io_next_1(rptr_io_next_1),
    .io_enable_0(rptr_io_enable_0),
    .io_enable_1(rptr_io_enable_1),
    .io_done_0(rptr_io_done_0),
    .io_config_chain_0(rptr_io_config_chain_0)
  );
  SRAM_10 mems_0_0 (
    .clock(mems_0_0_clock),
    .reset(mems_0_0_reset),
    .io_raddr(mems_0_0_io_raddr),
    .io_wen(mems_0_0_io_wen),
    .io_waddr(mems_0_0_io_waddr),
    .io_wdata_addr(mems_0_0_io_wdata_addr),
    .io_wdata_isWr(mems_0_0_io_wdata_isWr),
    .io_wdata_size(mems_0_0_io_wdata_size),
    .io_rdata_addr(mems_0_0_io_rdata_addr),
    .io_rdata_isWr(mems_0_0_io_rdata_isWr),
    .io_rdata_size(mems_0_0_io_rdata_size)
  );
  MuxN_2 MuxN (
    .io_ins_0_addr(MuxN_io_ins_0_addr),
    .io_ins_0_isWr(MuxN_io_ins_0_isWr),
    .io_ins_0_size(MuxN_io_ins_0_size),
    .io_out_addr(MuxN_io_out_addr),
    .io_out_isWr(MuxN_io_out_isWr),
    .io_out_size(MuxN_io_out_size)
  );
  assign _T_21 = 9'h100 - sizeUDC_io_out;
  assign _T_22 = $unsigned(_T_21);
  assign remainingSlots = _T_22[8:0];
  assign empty = sizeUDC_io_out < 9'h1;
  assign almostEmpty = sizeUDC_io_nextDec < 9'h1;
  assign full = remainingSlots < 9'h1;
  assign _T_34 = ~ full;
  assign writeEn = io_enqVld & _T_34;
  assign _T_35 = ~ empty;
  assign readEn = io_deqVld & _T_35;
  assign nextHeadLocalAddr = rptr_io_done_0 ? rptr_io_next_1 : rptr_io_out_1;
  assign _T_79 = readEn ? nextHeadLocalAddr : rptr_io_out_1;
  assign _T_81 = wptr_io_out_0 == 9'h0;
  assign _T_82 = writeEn & _T_81;
  assign io_deq_0_addr = MuxN_io_out_addr;
  assign io_deq_0_isWr = MuxN_io_out_isWr;
  assign io_deq_0_size = MuxN_io_out_size;
  assign io_full = full;
  assign io_empty = empty;
  assign io_almostEmpty = almostEmpty;
  assign sizeUDC_io_strideInc = 9'h1;
  assign sizeUDC_io_strideDec = 9'h1;
  assign sizeUDC_io_inc = writeEn;
  assign sizeUDC_io_dec = readEn;
  assign sizeUDC_clock = clock;
  assign sizeUDC_reset = reset;
  assign wptr_io_enable_0 = writeEn;
  assign wptr_io_enable_1 = writeEn;
  assign wptr_io_config_chain_0 = 1'h1;
  assign wptr_clock = clock;
  assign wptr_reset = reset;
  assign rptr_io_enable_0 = readEn;
  assign rptr_io_enable_1 = readEn;
  assign rptr_io_config_chain_0 = 1'h1;
  assign rptr_clock = clock;
  assign rptr_reset = reset;
  assign mems_0_0_io_raddr = _T_79[7:0];
  assign mems_0_0_io_wen = _T_82;
  assign mems_0_0_io_waddr = wptr_io_out_1[7:0];
  assign mems_0_0_io_wdata_addr = wdata_0_addr;
  assign mems_0_0_io_wdata_isWr = wdata_0_isWr;
  assign mems_0_0_io_wdata_size = wdata_0_size;
  assign mems_0_0_clock = clock;
  assign mems_0_0_reset = reset;
  assign wdata_0_addr = io_enq_0_addr;
  assign wdata_0_isWr = io_enq_0_isWr;
  assign wdata_0_size = io_enq_0_size;
  assign MuxN_io_ins_0_addr = mems_0_0_io_rdata_addr;
  assign MuxN_io_ins_0_isWr = mems_0_0_io_rdata_isWr;
  assign MuxN_io_ins_0_size = mems_0_0_io_rdata_size;
endmodule
module RetimeWrapper_579(
  input         clock,
  input         reset,
  input  [63:0] io_in,
  output [63:0] io_out
);
  wire [63:0] sr_out;
  wire [63:0] sr_in;
  wire  sr_flow;
  wire  sr_reset;
  wire  sr_clock;
  RetimeShiftRegister #(.WIDTH(64), .STAGES(1)) sr (
    .out(sr_out),
    .in(sr_in),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out;
  assign sr_in = io_in;
  assign sr_flow = 1'h1;
  assign sr_reset = reset;
  assign sr_clock = clock;
endmodule
module FF_136(
  input         clock,
  input         reset,
  input  [63:0] io_in,
  input  [63:0] io_init,
  input         io_reset,
  output [63:0] io_out,
  input         io_enable
);
  wire [63:0] d;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire [63:0] RetimeWrapper_io_in;
  wire [63:0] RetimeWrapper_io_out;
  wire [63:0] _T_11;
  wire [63:0] _GEN_0;
  wire [63:0] _GEN_1;
  RetimeWrapper_579 RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _GEN_0 = io_reset ? io_init : _T_11;
  assign _GEN_1 = io_enable ? io_in : _GEN_0;
  assign io_out = _T_11;
  assign d = _GEN_1;
  assign RetimeWrapper_io_in = d;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_11 = RetimeWrapper_io_out;
endmodule
module RetimeWrapper_580(
  input         clock,
  input         reset,
  input  [15:0] io_in,
  output [15:0] io_out
);
  wire [15:0] sr_out;
  wire [15:0] sr_in;
  wire  sr_flow;
  wire  sr_reset;
  wire  sr_clock;
  RetimeShiftRegister #(.WIDTH(16), .STAGES(1)) sr (
    .out(sr_out),
    .in(sr_in),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out;
  assign sr_in = io_in;
  assign sr_flow = 1'h1;
  assign sr_reset = reset;
  assign sr_clock = clock;
endmodule
module FF_137(
  input         clock,
  input         reset,
  input  [15:0] io_in,
  output [15:0] io_out,
  input         io_enable
);
  wire [15:0] d;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire [15:0] RetimeWrapper_io_in;
  wire [15:0] RetimeWrapper_io_out;
  wire [15:0] _T_11;
  wire [15:0] _GEN_1;
  RetimeWrapper_580 RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _GEN_1 = io_enable ? io_in : _T_11;
  assign io_out = _T_11;
  assign d = _GEN_1;
  assign RetimeWrapper_io_in = d;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_11 = RetimeWrapper_io_out;
endmodule
module Counter_15(
  input         clock,
  input         reset,
  input  [15:0] io_max,
  input  [15:0] io_stride,
  output [15:0] io_out,
  output        io_last,
  input         io_reset,
  input         io_enable,
  output        io_done
);
  wire  reg$_clock;
  wire  reg$_reset;
  wire [15:0] reg$_io_in;
  wire [15:0] reg$_io_out;
  wire  reg$_io_enable;
  wire  _T_11;
  wire [16:0] count;
  wire [16:0] _GEN_1;
  wire [17:0] _T_13;
  wire [16:0] newval;
  wire [16:0] _GEN_2;
  wire  isMax;
  wire [16:0] next;
  wire [16:0] _GEN_0;
  wire  _T_15;
  FF_137 reg$ (
    .clock(reg$_clock),
    .reset(reg$_reset),
    .io_in(reg$_io_in),
    .io_out(reg$_io_out),
    .io_enable(reg$_io_enable)
  );
  assign _T_11 = io_reset | io_enable;
  assign count = {1'h0,reg$_io_out};
  assign _GEN_1 = {{1'd0}, io_stride};
  assign _T_13 = count + _GEN_1;
  assign newval = _T_13[16:0];
  assign _GEN_2 = {{1'd0}, io_max};
  assign isMax = newval >= _GEN_2;
  assign next = isMax ? 17'h0 : newval;
  assign _GEN_0 = io_reset ? 17'h0 : next;
  assign _T_15 = io_enable & isMax;
  assign io_out = count[15:0];
  assign io_last = isMax;
  assign io_done = _T_15;
  assign reg$_io_in = _GEN_0[15:0];
  assign reg$_io_enable = _T_11;
  assign reg$_clock = clock;
  assign reg$_reset = reset;
endmodule
module MuxN_4(
  input   io_ins_0,
  input   io_ins_1,
  input   io_sel,
  output  io_out
);
  wire  _GEN_0;
  wire  _GEN_1;
  assign _GEN_1 = io_sel ? io_ins_1 : io_ins_0;
  assign io_out = _GEN_0;
  assign _GEN_0 = _GEN_1;
endmodule
module RetimeWrapper_582(
  input        clock,
  input        reset,
  input  [9:0] io_in,
  output [9:0] io_out
);
  wire [9:0] sr_out;
  wire [9:0] sr_in;
  wire  sr_flow;
  wire  sr_reset;
  wire  sr_clock;
  RetimeShiftRegister #(.WIDTH(10), .STAGES(1)) sr (
    .out(sr_out),
    .in(sr_in),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out;
  assign sr_in = io_in;
  assign sr_flow = 1'h1;
  assign sr_reset = reset;
  assign sr_clock = clock;
endmodule
module FF_139(
  input        clock,
  input        reset,
  input  [9:0] io_in,
  output [9:0] io_out,
  input        io_enable
);
  wire [9:0] d;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire [9:0] RetimeWrapper_io_in;
  wire [9:0] RetimeWrapper_io_out;
  wire [9:0] _T_11;
  wire [9:0] _GEN_1;
  RetimeWrapper_582 RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _GEN_1 = io_enable ? io_in : _T_11;
  assign io_out = _T_11;
  assign d = _GEN_1;
  assign RetimeWrapper_io_in = d;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_11 = RetimeWrapper_io_out;
endmodule
module Counter_17(
  input        clock,
  input        reset,
  output [9:0] io_out,
  input        io_reset,
  input        io_enable
);
  wire  reg$_clock;
  wire  reg$_reset;
  wire [9:0] reg$_io_in;
  wire [9:0] reg$_io_out;
  wire  reg$_io_enable;
  wire  _T_11;
  wire [10:0] count;
  wire [11:0] _T_13;
  wire [10:0] newval;
  wire  isMax;
  wire [10:0] next;
  wire [10:0] _GEN_0;
  FF_139 reg$ (
    .clock(reg$_clock),
    .reset(reg$_reset),
    .io_in(reg$_io_in),
    .io_out(reg$_io_out),
    .io_enable(reg$_io_enable)
  );
  assign _T_11 = io_reset | io_enable;
  assign count = {1'h0,reg$_io_out};
  assign _T_13 = count + 11'h1;
  assign newval = _T_13[10:0];
  assign isMax = newval >= 11'h3ff;
  assign next = isMax ? 11'h0 : newval;
  assign _GEN_0 = io_reset ? 11'h0 : next;
  assign io_out = count[9:0];
  assign reg$_io_in = _GEN_0[9:0];
  assign reg$_io_enable = _T_11;
  assign reg$_clock = clock;
  assign reg$_reset = reset;
endmodule
module MuxN_5(
  input   io_ins_0,
  output  io_out
);
  assign io_out = io_ins_0;
endmodule
module MuxN_6(
  input         io_ins_0_valid,
  input  [31:0] io_ins_0_bits_wdata_0,
  input  [31:0] io_ins_0_bits_wdata_1,
  input  [31:0] io_ins_0_bits_wdata_2,
  input  [31:0] io_ins_0_bits_wdata_3,
  input  [31:0] io_ins_0_bits_wdata_4,
  input  [31:0] io_ins_0_bits_wdata_5,
  input  [31:0] io_ins_0_bits_wdata_6,
  input  [31:0] io_ins_0_bits_wdata_7,
  input  [31:0] io_ins_0_bits_wdata_8,
  input  [31:0] io_ins_0_bits_wdata_9,
  input  [31:0] io_ins_0_bits_wdata_10,
  input  [31:0] io_ins_0_bits_wdata_11,
  input  [31:0] io_ins_0_bits_wdata_12,
  input  [31:0] io_ins_0_bits_wdata_13,
  input  [31:0] io_ins_0_bits_wdata_14,
  input  [31:0] io_ins_0_bits_wdata_15,
  input         io_ins_0_bits_wstrb_0,
  input         io_ins_0_bits_wstrb_1,
  input         io_ins_0_bits_wstrb_2,
  input         io_ins_0_bits_wstrb_3,
  input         io_ins_0_bits_wstrb_4,
  input         io_ins_0_bits_wstrb_5,
  input         io_ins_0_bits_wstrb_6,
  input         io_ins_0_bits_wstrb_7,
  input         io_ins_0_bits_wstrb_8,
  input         io_ins_0_bits_wstrb_9,
  input         io_ins_0_bits_wstrb_10,
  input         io_ins_0_bits_wstrb_11,
  input         io_ins_0_bits_wstrb_12,
  input         io_ins_0_bits_wstrb_13,
  input         io_ins_0_bits_wstrb_14,
  input         io_ins_0_bits_wstrb_15,
  input         io_ins_0_bits_wstrb_16,
  input         io_ins_0_bits_wstrb_17,
  input         io_ins_0_bits_wstrb_18,
  input         io_ins_0_bits_wstrb_19,
  input         io_ins_0_bits_wstrb_20,
  input         io_ins_0_bits_wstrb_21,
  input         io_ins_0_bits_wstrb_22,
  input         io_ins_0_bits_wstrb_23,
  input         io_ins_0_bits_wstrb_24,
  input         io_ins_0_bits_wstrb_25,
  input         io_ins_0_bits_wstrb_26,
  input         io_ins_0_bits_wstrb_27,
  input         io_ins_0_bits_wstrb_28,
  input         io_ins_0_bits_wstrb_29,
  input         io_ins_0_bits_wstrb_30,
  input         io_ins_0_bits_wstrb_31,
  input         io_ins_0_bits_wstrb_32,
  input         io_ins_0_bits_wstrb_33,
  input         io_ins_0_bits_wstrb_34,
  input         io_ins_0_bits_wstrb_35,
  input         io_ins_0_bits_wstrb_36,
  input         io_ins_0_bits_wstrb_37,
  input         io_ins_0_bits_wstrb_38,
  input         io_ins_0_bits_wstrb_39,
  input         io_ins_0_bits_wstrb_40,
  input         io_ins_0_bits_wstrb_41,
  input         io_ins_0_bits_wstrb_42,
  input         io_ins_0_bits_wstrb_43,
  input         io_ins_0_bits_wstrb_44,
  input         io_ins_0_bits_wstrb_45,
  input         io_ins_0_bits_wstrb_46,
  input         io_ins_0_bits_wstrb_47,
  input         io_ins_0_bits_wstrb_48,
  input         io_ins_0_bits_wstrb_49,
  input         io_ins_0_bits_wstrb_50,
  input         io_ins_0_bits_wstrb_51,
  input         io_ins_0_bits_wstrb_52,
  input         io_ins_0_bits_wstrb_53,
  input         io_ins_0_bits_wstrb_54,
  input         io_ins_0_bits_wstrb_55,
  input         io_ins_0_bits_wstrb_56,
  input         io_ins_0_bits_wstrb_57,
  input         io_ins_0_bits_wstrb_58,
  input         io_ins_0_bits_wstrb_59,
  input         io_ins_0_bits_wstrb_60,
  input         io_ins_0_bits_wstrb_61,
  input         io_ins_0_bits_wstrb_62,
  input         io_ins_0_bits_wstrb_63,
  output        io_out_valid,
  output [31:0] io_out_bits_wdata_0,
  output [31:0] io_out_bits_wdata_1,
  output [31:0] io_out_bits_wdata_2,
  output [31:0] io_out_bits_wdata_3,
  output [31:0] io_out_bits_wdata_4,
  output [31:0] io_out_bits_wdata_5,
  output [31:0] io_out_bits_wdata_6,
  output [31:0] io_out_bits_wdata_7,
  output [31:0] io_out_bits_wdata_8,
  output [31:0] io_out_bits_wdata_9,
  output [31:0] io_out_bits_wdata_10,
  output [31:0] io_out_bits_wdata_11,
  output [31:0] io_out_bits_wdata_12,
  output [31:0] io_out_bits_wdata_13,
  output [31:0] io_out_bits_wdata_14,
  output [31:0] io_out_bits_wdata_15,
  output        io_out_bits_wstrb_0,
  output        io_out_bits_wstrb_1,
  output        io_out_bits_wstrb_2,
  output        io_out_bits_wstrb_3,
  output        io_out_bits_wstrb_4,
  output        io_out_bits_wstrb_5,
  output        io_out_bits_wstrb_6,
  output        io_out_bits_wstrb_7,
  output        io_out_bits_wstrb_8,
  output        io_out_bits_wstrb_9,
  output        io_out_bits_wstrb_10,
  output        io_out_bits_wstrb_11,
  output        io_out_bits_wstrb_12,
  output        io_out_bits_wstrb_13,
  output        io_out_bits_wstrb_14,
  output        io_out_bits_wstrb_15,
  output        io_out_bits_wstrb_16,
  output        io_out_bits_wstrb_17,
  output        io_out_bits_wstrb_18,
  output        io_out_bits_wstrb_19,
  output        io_out_bits_wstrb_20,
  output        io_out_bits_wstrb_21,
  output        io_out_bits_wstrb_22,
  output        io_out_bits_wstrb_23,
  output        io_out_bits_wstrb_24,
  output        io_out_bits_wstrb_25,
  output        io_out_bits_wstrb_26,
  output        io_out_bits_wstrb_27,
  output        io_out_bits_wstrb_28,
  output        io_out_bits_wstrb_29,
  output        io_out_bits_wstrb_30,
  output        io_out_bits_wstrb_31,
  output        io_out_bits_wstrb_32,
  output        io_out_bits_wstrb_33,
  output        io_out_bits_wstrb_34,
  output        io_out_bits_wstrb_35,
  output        io_out_bits_wstrb_36,
  output        io_out_bits_wstrb_37,
  output        io_out_bits_wstrb_38,
  output        io_out_bits_wstrb_39,
  output        io_out_bits_wstrb_40,
  output        io_out_bits_wstrb_41,
  output        io_out_bits_wstrb_42,
  output        io_out_bits_wstrb_43,
  output        io_out_bits_wstrb_44,
  output        io_out_bits_wstrb_45,
  output        io_out_bits_wstrb_46,
  output        io_out_bits_wstrb_47,
  output        io_out_bits_wstrb_48,
  output        io_out_bits_wstrb_49,
  output        io_out_bits_wstrb_50,
  output        io_out_bits_wstrb_51,
  output        io_out_bits_wstrb_52,
  output        io_out_bits_wstrb_53,
  output        io_out_bits_wstrb_54,
  output        io_out_bits_wstrb_55,
  output        io_out_bits_wstrb_56,
  output        io_out_bits_wstrb_57,
  output        io_out_bits_wstrb_58,
  output        io_out_bits_wstrb_59,
  output        io_out_bits_wstrb_60,
  output        io_out_bits_wstrb_61,
  output        io_out_bits_wstrb_62,
  output        io_out_bits_wstrb_63
);
  assign io_out_valid = io_ins_0_valid;
  assign io_out_bits_wdata_0 = io_ins_0_bits_wdata_0;
  assign io_out_bits_wdata_1 = io_ins_0_bits_wdata_1;
  assign io_out_bits_wdata_2 = io_ins_0_bits_wdata_2;
  assign io_out_bits_wdata_3 = io_ins_0_bits_wdata_3;
  assign io_out_bits_wdata_4 = io_ins_0_bits_wdata_4;
  assign io_out_bits_wdata_5 = io_ins_0_bits_wdata_5;
  assign io_out_bits_wdata_6 = io_ins_0_bits_wdata_6;
  assign io_out_bits_wdata_7 = io_ins_0_bits_wdata_7;
  assign io_out_bits_wdata_8 = io_ins_0_bits_wdata_8;
  assign io_out_bits_wdata_9 = io_ins_0_bits_wdata_9;
  assign io_out_bits_wdata_10 = io_ins_0_bits_wdata_10;
  assign io_out_bits_wdata_11 = io_ins_0_bits_wdata_11;
  assign io_out_bits_wdata_12 = io_ins_0_bits_wdata_12;
  assign io_out_bits_wdata_13 = io_ins_0_bits_wdata_13;
  assign io_out_bits_wdata_14 = io_ins_0_bits_wdata_14;
  assign io_out_bits_wdata_15 = io_ins_0_bits_wdata_15;
  assign io_out_bits_wstrb_0 = io_ins_0_bits_wstrb_0;
  assign io_out_bits_wstrb_1 = io_ins_0_bits_wstrb_1;
  assign io_out_bits_wstrb_2 = io_ins_0_bits_wstrb_2;
  assign io_out_bits_wstrb_3 = io_ins_0_bits_wstrb_3;
  assign io_out_bits_wstrb_4 = io_ins_0_bits_wstrb_4;
  assign io_out_bits_wstrb_5 = io_ins_0_bits_wstrb_5;
  assign io_out_bits_wstrb_6 = io_ins_0_bits_wstrb_6;
  assign io_out_bits_wstrb_7 = io_ins_0_bits_wstrb_7;
  assign io_out_bits_wstrb_8 = io_ins_0_bits_wstrb_8;
  assign io_out_bits_wstrb_9 = io_ins_0_bits_wstrb_9;
  assign io_out_bits_wstrb_10 = io_ins_0_bits_wstrb_10;
  assign io_out_bits_wstrb_11 = io_ins_0_bits_wstrb_11;
  assign io_out_bits_wstrb_12 = io_ins_0_bits_wstrb_12;
  assign io_out_bits_wstrb_13 = io_ins_0_bits_wstrb_13;
  assign io_out_bits_wstrb_14 = io_ins_0_bits_wstrb_14;
  assign io_out_bits_wstrb_15 = io_ins_0_bits_wstrb_15;
  assign io_out_bits_wstrb_16 = io_ins_0_bits_wstrb_16;
  assign io_out_bits_wstrb_17 = io_ins_0_bits_wstrb_17;
  assign io_out_bits_wstrb_18 = io_ins_0_bits_wstrb_18;
  assign io_out_bits_wstrb_19 = io_ins_0_bits_wstrb_19;
  assign io_out_bits_wstrb_20 = io_ins_0_bits_wstrb_20;
  assign io_out_bits_wstrb_21 = io_ins_0_bits_wstrb_21;
  assign io_out_bits_wstrb_22 = io_ins_0_bits_wstrb_22;
  assign io_out_bits_wstrb_23 = io_ins_0_bits_wstrb_23;
  assign io_out_bits_wstrb_24 = io_ins_0_bits_wstrb_24;
  assign io_out_bits_wstrb_25 = io_ins_0_bits_wstrb_25;
  assign io_out_bits_wstrb_26 = io_ins_0_bits_wstrb_26;
  assign io_out_bits_wstrb_27 = io_ins_0_bits_wstrb_27;
  assign io_out_bits_wstrb_28 = io_ins_0_bits_wstrb_28;
  assign io_out_bits_wstrb_29 = io_ins_0_bits_wstrb_29;
  assign io_out_bits_wstrb_30 = io_ins_0_bits_wstrb_30;
  assign io_out_bits_wstrb_31 = io_ins_0_bits_wstrb_31;
  assign io_out_bits_wstrb_32 = io_ins_0_bits_wstrb_32;
  assign io_out_bits_wstrb_33 = io_ins_0_bits_wstrb_33;
  assign io_out_bits_wstrb_34 = io_ins_0_bits_wstrb_34;
  assign io_out_bits_wstrb_35 = io_ins_0_bits_wstrb_35;
  assign io_out_bits_wstrb_36 = io_ins_0_bits_wstrb_36;
  assign io_out_bits_wstrb_37 = io_ins_0_bits_wstrb_37;
  assign io_out_bits_wstrb_38 = io_ins_0_bits_wstrb_38;
  assign io_out_bits_wstrb_39 = io_ins_0_bits_wstrb_39;
  assign io_out_bits_wstrb_40 = io_ins_0_bits_wstrb_40;
  assign io_out_bits_wstrb_41 = io_ins_0_bits_wstrb_41;
  assign io_out_bits_wstrb_42 = io_ins_0_bits_wstrb_42;
  assign io_out_bits_wstrb_43 = io_ins_0_bits_wstrb_43;
  assign io_out_bits_wstrb_44 = io_ins_0_bits_wstrb_44;
  assign io_out_bits_wstrb_45 = io_ins_0_bits_wstrb_45;
  assign io_out_bits_wstrb_46 = io_ins_0_bits_wstrb_46;
  assign io_out_bits_wstrb_47 = io_ins_0_bits_wstrb_47;
  assign io_out_bits_wstrb_48 = io_ins_0_bits_wstrb_48;
  assign io_out_bits_wstrb_49 = io_ins_0_bits_wstrb_49;
  assign io_out_bits_wstrb_50 = io_ins_0_bits_wstrb_50;
  assign io_out_bits_wstrb_51 = io_ins_0_bits_wstrb_51;
  assign io_out_bits_wstrb_52 = io_ins_0_bits_wstrb_52;
  assign io_out_bits_wstrb_53 = io_ins_0_bits_wstrb_53;
  assign io_out_bits_wstrb_54 = io_ins_0_bits_wstrb_54;
  assign io_out_bits_wstrb_55 = io_ins_0_bits_wstrb_55;
  assign io_out_bits_wstrb_56 = io_ins_0_bits_wstrb_56;
  assign io_out_bits_wstrb_57 = io_ins_0_bits_wstrb_57;
  assign io_out_bits_wstrb_58 = io_ins_0_bits_wstrb_58;
  assign io_out_bits_wstrb_59 = io_ins_0_bits_wstrb_59;
  assign io_out_bits_wstrb_60 = io_ins_0_bits_wstrb_60;
  assign io_out_bits_wstrb_61 = io_ins_0_bits_wstrb_61;
  assign io_out_bits_wstrb_62 = io_ins_0_bits_wstrb_62;
  assign io_out_bits_wstrb_63 = io_ins_0_bits_wstrb_63;
endmodule
module MuxN_8(
  input         io_ins_0_valid,
  input  [63:0] io_ins_0_bits_addr,
  input  [31:0] io_ins_0_bits_size,
  input         io_ins_0_bits_isWr,
  input  [25:0] io_ins_0_bits_tag_uid,
  input  [5:0]  io_ins_0_bits_tag_streamId,
  input         io_ins_1_valid,
  input  [63:0] io_ins_1_bits_addr,
  input  [31:0] io_ins_1_bits_size,
  input         io_ins_1_bits_isWr,
  input  [25:0] io_ins_1_bits_tag_uid,
  input  [5:0]  io_ins_1_bits_tag_streamId,
  input         io_sel,
  output        io_out_valid,
  output [63:0] io_out_bits_addr,
  output [31:0] io_out_bits_size,
  output        io_out_bits_isWr,
  output [25:0] io_out_bits_tag_uid,
  output [5:0]  io_out_bits_tag_streamId
);
  wire  _GEN_8;
  wire [63:0] _GEN_9;
  wire [31:0] _GEN_10;
  wire  _GEN_12;
  wire [25:0] _GEN_13;
  wire [5:0] _GEN_14;
  wire [5:0] _GEN_1_bits_tag_streamId;
  wire [25:0] _GEN_2_bits_tag_uid;
  wire  _GEN_3_bits_isWr;
  wire [31:0] _GEN_5_bits_size;
  wire [63:0] _GEN_6_bits_addr;
  wire  _GEN_7_valid;
  assign _GEN_8 = io_sel ? io_ins_1_valid : io_ins_0_valid;
  assign _GEN_9 = io_sel ? io_ins_1_bits_addr : io_ins_0_bits_addr;
  assign _GEN_10 = io_sel ? io_ins_1_bits_size : io_ins_0_bits_size;
  assign _GEN_12 = io_sel ? io_ins_1_bits_isWr : io_ins_0_bits_isWr;
  assign _GEN_13 = io_sel ? io_ins_1_bits_tag_uid : io_ins_0_bits_tag_uid;
  assign _GEN_14 = io_sel ? io_ins_1_bits_tag_streamId : io_ins_0_bits_tag_streamId;
  assign io_out_valid = _GEN_7_valid;
  assign io_out_bits_addr = _GEN_6_bits_addr;
  assign io_out_bits_size = _GEN_5_bits_size;
  assign io_out_bits_isWr = _GEN_3_bits_isWr;
  assign io_out_bits_tag_uid = _GEN_2_bits_tag_uid;
  assign io_out_bits_tag_streamId = _GEN_1_bits_tag_streamId;
  assign _GEN_1_bits_tag_streamId = _GEN_14;
  assign _GEN_2_bits_tag_uid = _GEN_13;
  assign _GEN_3_bits_isWr = _GEN_12;
  assign _GEN_5_bits_size = _GEN_10;
  assign _GEN_6_bits_addr = _GEN_9;
  assign _GEN_7_valid = _GEN_8;
endmodule
module RetimeWrapper_586(
  input        clock,
  input        reset,
  input  [5:0] io_in,
  output [5:0] io_out
);
  wire [5:0] sr_out;
  wire [5:0] sr_in;
  wire  sr_flow;
  wire  sr_reset;
  wire  sr_clock;
  RetimeShiftRegister #(.WIDTH(6), .STAGES(1)) sr (
    .out(sr_out),
    .in(sr_in),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out;
  assign sr_in = io_in;
  assign sr_flow = 1'h1;
  assign sr_reset = reset;
  assign sr_clock = clock;
endmodule
module FF_143(
  input        clock,
  input        reset,
  input  [5:0] io_in,
  output [5:0] io_out,
  input        io_enable
);
  wire [5:0] d;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire [5:0] RetimeWrapper_io_in;
  wire [5:0] RetimeWrapper_io_out;
  wire [5:0] _T_11;
  wire [5:0] _GEN_1;
  RetimeWrapper_586 RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _GEN_1 = io_enable ? io_in : _T_11;
  assign io_out = _T_11;
  assign d = _GEN_1;
  assign RetimeWrapper_io_in = d;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_11 = RetimeWrapper_io_out;
endmodule
module FF_145(
  input         clock,
  input         reset,
  input  [31:0] io_in,
  output [31:0] io_out,
  input         io_enable
);
  wire [31:0] d;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire [31:0] RetimeWrapper_io_in;
  wire [31:0] RetimeWrapper_io_out;
  wire [31:0] _T_11;
  wire [31:0] _GEN_1;
  RetimeWrapper_6 RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _GEN_1 = io_enable ? io_in : _T_11;
  assign io_out = _T_11;
  assign d = _GEN_1;
  assign RetimeWrapper_io_in = d;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_11 = RetimeWrapper_io_out;
endmodule
module Counter_18(
  input         clock,
  input         reset,
  output [63:0] io_out,
  input         io_reset,
  input         io_enable
);
  wire  reg$_clock;
  wire  reg$_reset;
  wire [63:0] reg$_io_in;
  wire [63:0] reg$_io_init;
  wire  reg$_io_reset;
  wire [63:0] reg$_io_out;
  wire  reg$_io_enable;
  wire  _T_11;
  wire [64:0] count;
  wire [65:0] _T_13;
  wire [64:0] newval;
  wire  isMax;
  wire [64:0] next;
  wire [64:0] _GEN_0;
  FF_136 reg$ (
    .clock(reg$_clock),
    .reset(reg$_reset),
    .io_in(reg$_io_in),
    .io_init(reg$_io_init),
    .io_reset(reg$_io_reset),
    .io_out(reg$_io_out),
    .io_enable(reg$_io_enable)
  );
  assign _T_11 = io_reset | io_enable;
  assign count = {1'h0,reg$_io_out};
  assign _T_13 = count + 65'h1;
  assign newval = _T_13[64:0];
  assign isMax = newval >= 65'hffffffff;
  assign next = isMax ? 65'h0 : newval;
  assign _GEN_0 = io_reset ? 65'h0 : next;
  assign io_out = count[63:0];
  assign reg$_io_in = _GEN_0[63:0];
  assign reg$_io_init = 64'h0;
  assign reg$_io_reset = 1'h0;
  assign reg$_io_enable = _T_11;
  assign reg$_clock = clock;
  assign reg$_reset = reset;
endmodule
module RetimeWrapper_598(
  input        clock,
  input        reset,
  input  [4:0] io_in,
  output [4:0] io_out
);
  wire [4:0] sr_out;
  wire [4:0] sr_in;
  wire  sr_flow;
  wire  sr_reset;
  wire  sr_clock;
  RetimeShiftRegister #(.WIDTH(5), .STAGES(1)) sr (
    .out(sr_out),
    .in(sr_in),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out;
  assign sr_in = io_in;
  assign sr_flow = 1'h1;
  assign sr_reset = reset;
  assign sr_clock = clock;
endmodule
module FF_155(
  input        clock,
  input        reset,
  input  [4:0] io_in,
  output [4:0] io_out,
  input        io_enable
);
  wire [4:0] d;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire [4:0] RetimeWrapper_io_in;
  wire [4:0] RetimeWrapper_io_out;
  wire [4:0] _T_11;
  wire [4:0] _GEN_1;
  RetimeWrapper_598 RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _GEN_1 = io_enable ? io_in : _T_11;
  assign io_out = _T_11;
  assign d = _GEN_1;
  assign RetimeWrapper_io_in = d;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_11 = RetimeWrapper_io_out;
endmodule
module Counter_24(
  input        clock,
  input        reset,
  output [4:0] io_out,
  output [4:0] io_next,
  input        io_enable,
  output       io_done
);
  wire  reg$_clock;
  wire  reg$_reset;
  wire [4:0] reg$_io_in;
  wire [4:0] reg$_io_out;
  wire  reg$_io_enable;
  wire [5:0] count;
  wire [6:0] _T_13;
  wire [5:0] newval;
  wire  isMax;
  wire [5:0] next;
  wire  _T_15;
  FF_155 reg$ (
    .clock(reg$_clock),
    .reset(reg$_reset),
    .io_in(reg$_io_in),
    .io_out(reg$_io_out),
    .io_enable(reg$_io_enable)
  );
  assign count = {1'h0,reg$_io_out};
  assign _T_13 = count + 6'h1;
  assign newval = _T_13[5:0];
  assign isMax = newval >= 6'h10;
  assign next = isMax ? 6'h0 : newval;
  assign _T_15 = io_enable & isMax;
  assign io_out = count[4:0];
  assign io_next = next[4:0];
  assign io_done = _T_15;
  assign reg$_io_in = next[4:0];
  assign reg$_io_enable = io_enable;
  assign reg$_clock = clock;
  assign reg$_reset = reset;
endmodule
module CounterCore_8(
  input        clock,
  input        reset,
  output [4:0] io_out,
  output [4:0] io_next,
  input        io_enable,
  output       io_done
);
  wire  counter_clock;
  wire  counter_reset;
  wire [4:0] counter_io_out;
  wire [4:0] counter_io_next;
  wire  counter_io_enable;
  wire  counter_io_done;
  wire  depulser_clock;
  wire  depulser_reset;
  wire  depulser_io_in;
  wire  depulser_io_rst;
  wire  depulser_io_out;
  Counter_24 counter (
    .clock(counter_clock),
    .reset(counter_reset),
    .io_out(counter_io_out),
    .io_next(counter_io_next),
    .io_enable(counter_io_enable),
    .io_done(counter_io_done)
  );
  Depulser depulser (
    .clock(depulser_clock),
    .reset(depulser_reset),
    .io_in(depulser_io_in),
    .io_rst(depulser_io_rst),
    .io_out(depulser_io_out)
  );
  assign io_out = counter_io_out;
  assign io_next = counter_io_next;
  assign io_done = counter_io_done;
  assign counter_io_enable = io_enable;
  assign counter_clock = clock;
  assign counter_reset = reset;
  assign depulser_io_in = counter_io_done;
  assign depulser_io_rst = 1'h0;
  assign depulser_clock = clock;
  assign depulser_reset = reset;
endmodule
module CounterChainCore_4(
  input        clock,
  input        reset,
  output [4:0] io_out_0,
  output [4:0] io_out_1,
  output [4:0] io_next_0,
  output [4:0] io_next_1,
  input        io_enable_0,
  input        io_enable_1,
  output       io_done_0,
  input        io_config_chain_0
);
  wire  counters_0_clock;
  wire  counters_0_reset;
  wire [4:0] counters_0_io_out;
  wire [4:0] counters_0_io_next;
  wire  counters_0_io_enable;
  wire  counters_0_io_done;
  wire  counters_1_clock;
  wire  counters_1_reset;
  wire [4:0] counters_1_io_out;
  wire [4:0] counters_1_io_next;
  wire  counters_1_io_enable;
  wire  counters_1_io_done;
  wire  _T_69;
  CounterCore_8 counters_0 (
    .clock(counters_0_clock),
    .reset(counters_0_reset),
    .io_out(counters_0_io_out),
    .io_next(counters_0_io_next),
    .io_enable(counters_0_io_enable),
    .io_done(counters_0_io_done)
  );
  CounterCore_8 counters_1 (
    .clock(counters_1_clock),
    .reset(counters_1_reset),
    .io_out(counters_1_io_out),
    .io_next(counters_1_io_next),
    .io_enable(counters_1_io_enable),
    .io_done(counters_1_io_done)
  );
  assign _T_69 = io_config_chain_0 ? counters_0_io_done : io_enable_1;
  assign io_out_0 = counters_0_io_out;
  assign io_out_1 = counters_1_io_out;
  assign io_next_0 = counters_0_io_next;
  assign io_next_1 = counters_1_io_next;
  assign io_done_0 = counters_0_io_done;
  assign counters_0_io_enable = io_enable_0;
  assign counters_0_clock = clock;
  assign counters_0_reset = reset;
  assign counters_1_io_enable = _T_69;
  assign counters_1_clock = clock;
  assign counters_1_reset = reset;
endmodule
module SRAM_12(
  input         clock,
  input         reset,
  input  [3:0]  io_raddr,
  input         io_wen,
  input  [3:0]  io_waddr,
  input  [31:0] io_wdata,
  output [31:0] io_rdata
);
  wire [31:0] SRAMVerilogAWS_rdata;
  wire [31:0] SRAMVerilogAWS_wdata;
  wire  SRAMVerilogAWS_flow;
  wire  SRAMVerilogAWS_wen;
  wire  SRAMVerilogAWS_waddrEn;
  wire  SRAMVerilogAWS_raddrEn;
  wire [3:0] SRAMVerilogAWS_waddr;
  wire [3:0] SRAMVerilogAWS_raddr;
  wire  SRAMVerilogAWS_clk;
  wire  _T_8;
  wire  _T_9;
  reg  _T_12;
  reg [31:0] _RAND_0;
  reg [31:0] _T_15;
  reg [31:0] _RAND_1;
  wire [31:0] _T_16;
  wire [31:0] _T_18;
  SRAMVerilogAWS #(.DWIDTH(32), .WORDS(16), .AWIDTH(4)) SRAMVerilogAWS (
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .flow(SRAMVerilogAWS_flow),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_8 = io_raddr == io_waddr;
  assign _T_9 = io_wen & _T_8;
  assign _T_16 = _T_12 ? _T_15 : SRAMVerilogAWS_rdata;
  assign io_rdata = _T_18;
  assign SRAMVerilogAWS_wdata = io_wdata;
  assign SRAMVerilogAWS_flow = 1'h1;
  assign SRAMVerilogAWS_wen = io_wen;
  assign SRAMVerilogAWS_waddrEn = 1'h1;
  assign SRAMVerilogAWS_raddrEn = 1'h1;
  assign SRAMVerilogAWS_waddr = io_waddr;
  assign SRAMVerilogAWS_raddr = io_raddr;
  assign SRAMVerilogAWS_clk = clock;
  assign _T_18 = _T_16;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_12 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_15 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_12 <= 1'h0;
    end else begin
      _T_12 <= _T_9;
    end
    if (reset) begin
      _T_15 <= 32'h0;
    end else begin
      _T_15 <= io_wdata;
    end
  end
endmodule
module MuxN_16(
  input  [31:0] io_ins_0,
  input  [31:0] io_ins_1,
  input  [31:0] io_ins_2,
  input  [31:0] io_ins_3,
  input  [31:0] io_ins_4,
  input  [31:0] io_ins_5,
  input  [31:0] io_ins_6,
  input  [31:0] io_ins_7,
  input  [31:0] io_ins_8,
  input  [31:0] io_ins_9,
  input  [31:0] io_ins_10,
  input  [31:0] io_ins_11,
  input  [31:0] io_ins_12,
  input  [31:0] io_ins_13,
  input  [31:0] io_ins_14,
  input  [31:0] io_ins_15,
  input  [3:0]  io_sel,
  output [31:0] io_out
);
  wire [31:0] _GEN_0;
  wire [31:0] _GEN_1;
  wire [31:0] _GEN_2;
  wire [31:0] _GEN_3;
  wire [31:0] _GEN_4;
  wire [31:0] _GEN_5;
  wire [31:0] _GEN_6;
  wire [31:0] _GEN_7;
  wire [31:0] _GEN_8;
  wire [31:0] _GEN_9;
  wire [31:0] _GEN_10;
  wire [31:0] _GEN_11;
  wire [31:0] _GEN_12;
  wire [31:0] _GEN_13;
  wire [31:0] _GEN_14;
  wire [31:0] _GEN_15;
  assign _GEN_1 = 4'h1 == io_sel ? io_ins_1 : io_ins_0;
  assign _GEN_2 = 4'h2 == io_sel ? io_ins_2 : _GEN_1;
  assign _GEN_3 = 4'h3 == io_sel ? io_ins_3 : _GEN_2;
  assign _GEN_4 = 4'h4 == io_sel ? io_ins_4 : _GEN_3;
  assign _GEN_5 = 4'h5 == io_sel ? io_ins_5 : _GEN_4;
  assign _GEN_6 = 4'h6 == io_sel ? io_ins_6 : _GEN_5;
  assign _GEN_7 = 4'h7 == io_sel ? io_ins_7 : _GEN_6;
  assign _GEN_8 = 4'h8 == io_sel ? io_ins_8 : _GEN_7;
  assign _GEN_9 = 4'h9 == io_sel ? io_ins_9 : _GEN_8;
  assign _GEN_10 = 4'ha == io_sel ? io_ins_10 : _GEN_9;
  assign _GEN_11 = 4'hb == io_sel ? io_ins_11 : _GEN_10;
  assign _GEN_12 = 4'hc == io_sel ? io_ins_12 : _GEN_11;
  assign _GEN_13 = 4'hd == io_sel ? io_ins_13 : _GEN_12;
  assign _GEN_14 = 4'he == io_sel ? io_ins_14 : _GEN_13;
  assign _GEN_15 = 4'hf == io_sel ? io_ins_15 : _GEN_14;
  assign io_out = _GEN_0;
  assign _GEN_0 = _GEN_15;
endmodule
module FF_163(
  input        clock,
  input        reset,
  input  [3:0] io_in,
  output [3:0] io_out
);
  wire [3:0] d;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire [3:0] RetimeWrapper_io_in;
  wire [3:0] RetimeWrapper_io_out;
  wire [3:0] _T_11;
  RetimeWrapper_49 RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_out = _T_11;
  assign d = io_in;
  assign RetimeWrapper_io_in = d;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_11 = RetimeWrapper_io_out;
endmodule
module FIFOCore_2(
  input         clock,
  input         reset,
  input  [31:0] io_enq_0,
  input  [31:0] io_enq_1,
  input  [31:0] io_enq_2,
  input  [31:0] io_enq_3,
  input  [31:0] io_enq_4,
  input  [31:0] io_enq_5,
  input  [31:0] io_enq_6,
  input  [31:0] io_enq_7,
  input  [31:0] io_enq_8,
  input  [31:0] io_enq_9,
  input  [31:0] io_enq_10,
  input  [31:0] io_enq_11,
  input  [31:0] io_enq_12,
  input  [31:0] io_enq_13,
  input  [31:0] io_enq_14,
  input  [31:0] io_enq_15,
  input         io_enqVld,
  output [31:0] io_deq_0,
  output [31:0] io_deq_1,
  output [31:0] io_deq_2,
  output [31:0] io_deq_3,
  output [31:0] io_deq_4,
  output [31:0] io_deq_5,
  output [31:0] io_deq_6,
  output [31:0] io_deq_7,
  output [31:0] io_deq_8,
  output [31:0] io_deq_9,
  output [31:0] io_deq_10,
  output [31:0] io_deq_11,
  output [31:0] io_deq_12,
  output [31:0] io_deq_13,
  output [31:0] io_deq_14,
  output [31:0] io_deq_15,
  input         io_deqVld,
  output        io_full,
  output        io_empty,
  output        io_almostFull,
  output        io_almostEmpty,
  input         io_config_chainRead
);
  wire  sizeUDC_clock;
  wire  sizeUDC_reset;
  wire [8:0] sizeUDC_io_strideInc;
  wire [8:0] sizeUDC_io_strideDec;
  wire  sizeUDC_io_inc;
  wire  sizeUDC_io_dec;
  wire [8:0] sizeUDC_io_out;
  wire [8:0] sizeUDC_io_nextInc;
  wire [8:0] sizeUDC_io_nextDec;
  wire [9:0] _T_51;
  wire [9:0] _T_52;
  wire [8:0] remainingSlots;
  wire [9:0] _T_54;
  wire [9:0] _T_55;
  wire [8:0] nextRemainingSlots;
  wire [4:0] strideDec;
  wire [8:0] _GEN_0;
  wire  empty;
  wire  almostEmpty;
  wire  full;
  wire  almostFull;
  wire  _T_64;
  wire  writeEn;
  wire  _T_65;
  wire  readEn;
  wire  wptr_clock;
  wire  wptr_reset;
  wire [4:0] wptr_io_out_0;
  wire [4:0] wptr_io_out_1;
  wire [4:0] wptr_io_next_0;
  wire [4:0] wptr_io_next_1;
  wire  wptr_io_enable_0;
  wire  wptr_io_enable_1;
  wire  wptr_io_done_0;
  wire  wptr_io_config_chain_0;
  wire  rptrConfig_chain_0;
  wire  rptr_clock;
  wire  rptr_reset;
  wire [4:0] rptr_io_out_0;
  wire [4:0] rptr_io_out_1;
  wire [4:0] rptr_io_next_0;
  wire [4:0] rptr_io_next_1;
  wire  rptr_io_enable_0;
  wire  rptr_io_enable_1;
  wire  rptr_io_done_0;
  wire  rptr_io_config_chain_0;
  wire  _T_101;
  wire [4:0] _T_102;
  wire [4:0] nextHeadLocalAddr;
  wire  mems_0_0_clock;
  wire  mems_0_0_reset;
  wire [3:0] mems_0_0_io_raddr;
  wire  mems_0_0_io_wen;
  wire [3:0] mems_0_0_io_waddr;
  wire [31:0] mems_0_0_io_wdata;
  wire [31:0] mems_0_0_io_rdata;
  wire  mems_0_1_clock;
  wire  mems_0_1_reset;
  wire [3:0] mems_0_1_io_raddr;
  wire  mems_0_1_io_wen;
  wire [3:0] mems_0_1_io_waddr;
  wire [31:0] mems_0_1_io_wdata;
  wire [31:0] mems_0_1_io_rdata;
  wire  mems_0_2_clock;
  wire  mems_0_2_reset;
  wire [3:0] mems_0_2_io_raddr;
  wire  mems_0_2_io_wen;
  wire [3:0] mems_0_2_io_waddr;
  wire [31:0] mems_0_2_io_wdata;
  wire [31:0] mems_0_2_io_rdata;
  wire  mems_0_3_clock;
  wire  mems_0_3_reset;
  wire [3:0] mems_0_3_io_raddr;
  wire  mems_0_3_io_wen;
  wire [3:0] mems_0_3_io_waddr;
  wire [31:0] mems_0_3_io_wdata;
  wire [31:0] mems_0_3_io_rdata;
  wire  mems_0_4_clock;
  wire  mems_0_4_reset;
  wire [3:0] mems_0_4_io_raddr;
  wire  mems_0_4_io_wen;
  wire [3:0] mems_0_4_io_waddr;
  wire [31:0] mems_0_4_io_wdata;
  wire [31:0] mems_0_4_io_rdata;
  wire  mems_0_5_clock;
  wire  mems_0_5_reset;
  wire [3:0] mems_0_5_io_raddr;
  wire  mems_0_5_io_wen;
  wire [3:0] mems_0_5_io_waddr;
  wire [31:0] mems_0_5_io_wdata;
  wire [31:0] mems_0_5_io_rdata;
  wire  mems_0_6_clock;
  wire  mems_0_6_reset;
  wire [3:0] mems_0_6_io_raddr;
  wire  mems_0_6_io_wen;
  wire [3:0] mems_0_6_io_waddr;
  wire [31:0] mems_0_6_io_wdata;
  wire [31:0] mems_0_6_io_rdata;
  wire  mems_0_7_clock;
  wire  mems_0_7_reset;
  wire [3:0] mems_0_7_io_raddr;
  wire  mems_0_7_io_wen;
  wire [3:0] mems_0_7_io_waddr;
  wire [31:0] mems_0_7_io_wdata;
  wire [31:0] mems_0_7_io_rdata;
  wire  mems_0_8_clock;
  wire  mems_0_8_reset;
  wire [3:0] mems_0_8_io_raddr;
  wire  mems_0_8_io_wen;
  wire [3:0] mems_0_8_io_waddr;
  wire [31:0] mems_0_8_io_wdata;
  wire [31:0] mems_0_8_io_rdata;
  wire  mems_0_9_clock;
  wire  mems_0_9_reset;
  wire [3:0] mems_0_9_io_raddr;
  wire  mems_0_9_io_wen;
  wire [3:0] mems_0_9_io_waddr;
  wire [31:0] mems_0_9_io_wdata;
  wire [31:0] mems_0_9_io_rdata;
  wire  mems_0_10_clock;
  wire  mems_0_10_reset;
  wire [3:0] mems_0_10_io_raddr;
  wire  mems_0_10_io_wen;
  wire [3:0] mems_0_10_io_waddr;
  wire [31:0] mems_0_10_io_wdata;
  wire [31:0] mems_0_10_io_rdata;
  wire  mems_0_11_clock;
  wire  mems_0_11_reset;
  wire [3:0] mems_0_11_io_raddr;
  wire  mems_0_11_io_wen;
  wire [3:0] mems_0_11_io_waddr;
  wire [31:0] mems_0_11_io_wdata;
  wire [31:0] mems_0_11_io_rdata;
  wire  mems_0_12_clock;
  wire  mems_0_12_reset;
  wire [3:0] mems_0_12_io_raddr;
  wire  mems_0_12_io_wen;
  wire [3:0] mems_0_12_io_waddr;
  wire [31:0] mems_0_12_io_wdata;
  wire [31:0] mems_0_12_io_rdata;
  wire  mems_0_13_clock;
  wire  mems_0_13_reset;
  wire [3:0] mems_0_13_io_raddr;
  wire  mems_0_13_io_wen;
  wire [3:0] mems_0_13_io_waddr;
  wire [31:0] mems_0_13_io_wdata;
  wire [31:0] mems_0_13_io_rdata;
  wire  mems_0_14_clock;
  wire  mems_0_14_reset;
  wire [3:0] mems_0_14_io_raddr;
  wire  mems_0_14_io_wen;
  wire [3:0] mems_0_14_io_waddr;
  wire [31:0] mems_0_14_io_wdata;
  wire [31:0] mems_0_14_io_rdata;
  wire  mems_0_15_clock;
  wire  mems_0_15_reset;
  wire [3:0] mems_0_15_io_raddr;
  wire  mems_0_15_io_wen;
  wire [3:0] mems_0_15_io_waddr;
  wire [31:0] mems_0_15_io_wdata;
  wire [31:0] mems_0_15_io_rdata;
  wire [31:0] wdata_0;
  wire [31:0] wdata_1;
  wire [31:0] wdata_2;
  wire [31:0] wdata_3;
  wire [31:0] wdata_4;
  wire [31:0] wdata_5;
  wire [31:0] wdata_6;
  wire [31:0] wdata_7;
  wire [31:0] wdata_8;
  wire [31:0] wdata_9;
  wire [31:0] wdata_10;
  wire [31:0] wdata_11;
  wire [31:0] wdata_12;
  wire [31:0] wdata_13;
  wire [31:0] wdata_14;
  wire [31:0] wdata_15;
  wire [4:0] _T_154;
  wire [31:0] MuxN_io_ins_0;
  wire [31:0] MuxN_io_ins_1;
  wire [31:0] MuxN_io_ins_2;
  wire [31:0] MuxN_io_ins_3;
  wire [31:0] MuxN_io_ins_4;
  wire [31:0] MuxN_io_ins_5;
  wire [31:0] MuxN_io_ins_6;
  wire [31:0] MuxN_io_ins_7;
  wire [31:0] MuxN_io_ins_8;
  wire [31:0] MuxN_io_ins_9;
  wire [31:0] MuxN_io_ins_10;
  wire [31:0] MuxN_io_ins_11;
  wire [31:0] MuxN_io_ins_12;
  wire [31:0] MuxN_io_ins_13;
  wire [31:0] MuxN_io_ins_14;
  wire [31:0] MuxN_io_ins_15;
  wire [3:0] MuxN_io_sel;
  wire [31:0] MuxN_io_out;
  wire  FF_clock;
  wire  FF_reset;
  wire [3:0] FF_io_in;
  wire [3:0] FF_io_out;
  wire [4:0] _T_159;
  wire [3:0] _T_162;
  UpDownCtr sizeUDC (
    .clock(sizeUDC_clock),
    .reset(sizeUDC_reset),
    .io_strideInc(sizeUDC_io_strideInc),
    .io_strideDec(sizeUDC_io_strideDec),
    .io_inc(sizeUDC_io_inc),
    .io_dec(sizeUDC_io_dec),
    .io_out(sizeUDC_io_out),
    .io_nextInc(sizeUDC_io_nextInc),
    .io_nextDec(sizeUDC_io_nextDec)
  );
  CounterChainCore_4 wptr (
    .clock(wptr_clock),
    .reset(wptr_reset),
    .io_out_0(wptr_io_out_0),
    .io_out_1(wptr_io_out_1),
    .io_next_0(wptr_io_next_0),
    .io_next_1(wptr_io_next_1),
    .io_enable_0(wptr_io_enable_0),
    .io_enable_1(wptr_io_enable_1),
    .io_done_0(wptr_io_done_0),
    .io_config_chain_0(wptr_io_config_chain_0)
  );
  CounterChainCore_4 rptr (
    .clock(rptr_clock),
    .reset(rptr_reset),
    .io_out_0(rptr_io_out_0),
    .io_out_1(rptr_io_out_1),
    .io_next_0(rptr_io_next_0),
    .io_next_1(rptr_io_next_1),
    .io_enable_0(rptr_io_enable_0),
    .io_enable_1(rptr_io_enable_1),
    .io_done_0(rptr_io_done_0),
    .io_config_chain_0(rptr_io_config_chain_0)
  );
  SRAM_12 mems_0_0 (
    .clock(mems_0_0_clock),
    .reset(mems_0_0_reset),
    .io_raddr(mems_0_0_io_raddr),
    .io_wen(mems_0_0_io_wen),
    .io_waddr(mems_0_0_io_waddr),
    .io_wdata(mems_0_0_io_wdata),
    .io_rdata(mems_0_0_io_rdata)
  );
  SRAM_12 mems_0_1 (
    .clock(mems_0_1_clock),
    .reset(mems_0_1_reset),
    .io_raddr(mems_0_1_io_raddr),
    .io_wen(mems_0_1_io_wen),
    .io_waddr(mems_0_1_io_waddr),
    .io_wdata(mems_0_1_io_wdata),
    .io_rdata(mems_0_1_io_rdata)
  );
  SRAM_12 mems_0_2 (
    .clock(mems_0_2_clock),
    .reset(mems_0_2_reset),
    .io_raddr(mems_0_2_io_raddr),
    .io_wen(mems_0_2_io_wen),
    .io_waddr(mems_0_2_io_waddr),
    .io_wdata(mems_0_2_io_wdata),
    .io_rdata(mems_0_2_io_rdata)
  );
  SRAM_12 mems_0_3 (
    .clock(mems_0_3_clock),
    .reset(mems_0_3_reset),
    .io_raddr(mems_0_3_io_raddr),
    .io_wen(mems_0_3_io_wen),
    .io_waddr(mems_0_3_io_waddr),
    .io_wdata(mems_0_3_io_wdata),
    .io_rdata(mems_0_3_io_rdata)
  );
  SRAM_12 mems_0_4 (
    .clock(mems_0_4_clock),
    .reset(mems_0_4_reset),
    .io_raddr(mems_0_4_io_raddr),
    .io_wen(mems_0_4_io_wen),
    .io_waddr(mems_0_4_io_waddr),
    .io_wdata(mems_0_4_io_wdata),
    .io_rdata(mems_0_4_io_rdata)
  );
  SRAM_12 mems_0_5 (
    .clock(mems_0_5_clock),
    .reset(mems_0_5_reset),
    .io_raddr(mems_0_5_io_raddr),
    .io_wen(mems_0_5_io_wen),
    .io_waddr(mems_0_5_io_waddr),
    .io_wdata(mems_0_5_io_wdata),
    .io_rdata(mems_0_5_io_rdata)
  );
  SRAM_12 mems_0_6 (
    .clock(mems_0_6_clock),
    .reset(mems_0_6_reset),
    .io_raddr(mems_0_6_io_raddr),
    .io_wen(mems_0_6_io_wen),
    .io_waddr(mems_0_6_io_waddr),
    .io_wdata(mems_0_6_io_wdata),
    .io_rdata(mems_0_6_io_rdata)
  );
  SRAM_12 mems_0_7 (
    .clock(mems_0_7_clock),
    .reset(mems_0_7_reset),
    .io_raddr(mems_0_7_io_raddr),
    .io_wen(mems_0_7_io_wen),
    .io_waddr(mems_0_7_io_waddr),
    .io_wdata(mems_0_7_io_wdata),
    .io_rdata(mems_0_7_io_rdata)
  );
  SRAM_12 mems_0_8 (
    .clock(mems_0_8_clock),
    .reset(mems_0_8_reset),
    .io_raddr(mems_0_8_io_raddr),
    .io_wen(mems_0_8_io_wen),
    .io_waddr(mems_0_8_io_waddr),
    .io_wdata(mems_0_8_io_wdata),
    .io_rdata(mems_0_8_io_rdata)
  );
  SRAM_12 mems_0_9 (
    .clock(mems_0_9_clock),
    .reset(mems_0_9_reset),
    .io_raddr(mems_0_9_io_raddr),
    .io_wen(mems_0_9_io_wen),
    .io_waddr(mems_0_9_io_waddr),
    .io_wdata(mems_0_9_io_wdata),
    .io_rdata(mems_0_9_io_rdata)
  );
  SRAM_12 mems_0_10 (
    .clock(mems_0_10_clock),
    .reset(mems_0_10_reset),
    .io_raddr(mems_0_10_io_raddr),
    .io_wen(mems_0_10_io_wen),
    .io_waddr(mems_0_10_io_waddr),
    .io_wdata(mems_0_10_io_wdata),
    .io_rdata(mems_0_10_io_rdata)
  );
  SRAM_12 mems_0_11 (
    .clock(mems_0_11_clock),
    .reset(mems_0_11_reset),
    .io_raddr(mems_0_11_io_raddr),
    .io_wen(mems_0_11_io_wen),
    .io_waddr(mems_0_11_io_waddr),
    .io_wdata(mems_0_11_io_wdata),
    .io_rdata(mems_0_11_io_rdata)
  );
  SRAM_12 mems_0_12 (
    .clock(mems_0_12_clock),
    .reset(mems_0_12_reset),
    .io_raddr(mems_0_12_io_raddr),
    .io_wen(mems_0_12_io_wen),
    .io_waddr(mems_0_12_io_waddr),
    .io_wdata(mems_0_12_io_wdata),
    .io_rdata(mems_0_12_io_rdata)
  );
  SRAM_12 mems_0_13 (
    .clock(mems_0_13_clock),
    .reset(mems_0_13_reset),
    .io_raddr(mems_0_13_io_raddr),
    .io_wen(mems_0_13_io_wen),
    .io_waddr(mems_0_13_io_waddr),
    .io_wdata(mems_0_13_io_wdata),
    .io_rdata(mems_0_13_io_rdata)
  );
  SRAM_12 mems_0_14 (
    .clock(mems_0_14_clock),
    .reset(mems_0_14_reset),
    .io_raddr(mems_0_14_io_raddr),
    .io_wen(mems_0_14_io_wen),
    .io_waddr(mems_0_14_io_waddr),
    .io_wdata(mems_0_14_io_wdata),
    .io_rdata(mems_0_14_io_rdata)
  );
  SRAM_12 mems_0_15 (
    .clock(mems_0_15_clock),
    .reset(mems_0_15_reset),
    .io_raddr(mems_0_15_io_raddr),
    .io_wen(mems_0_15_io_wen),
    .io_waddr(mems_0_15_io_waddr),
    .io_wdata(mems_0_15_io_wdata),
    .io_rdata(mems_0_15_io_rdata)
  );
  MuxN_16 MuxN (
    .io_ins_0(MuxN_io_ins_0),
    .io_ins_1(MuxN_io_ins_1),
    .io_ins_2(MuxN_io_ins_2),
    .io_ins_3(MuxN_io_ins_3),
    .io_ins_4(MuxN_io_ins_4),
    .io_ins_5(MuxN_io_ins_5),
    .io_ins_6(MuxN_io_ins_6),
    .io_ins_7(MuxN_io_ins_7),
    .io_ins_8(MuxN_io_ins_8),
    .io_ins_9(MuxN_io_ins_9),
    .io_ins_10(MuxN_io_ins_10),
    .io_ins_11(MuxN_io_ins_11),
    .io_ins_12(MuxN_io_ins_12),
    .io_ins_13(MuxN_io_ins_13),
    .io_ins_14(MuxN_io_ins_14),
    .io_ins_15(MuxN_io_ins_15),
    .io_sel(MuxN_io_sel),
    .io_out(MuxN_io_out)
  );
  FF_163 FF (
    .clock(FF_clock),
    .reset(FF_reset),
    .io_in(FF_io_in),
    .io_out(FF_io_out)
  );
  assign _T_51 = 9'h100 - sizeUDC_io_out;
  assign _T_52 = $unsigned(_T_51);
  assign remainingSlots = _T_52[8:0];
  assign _T_54 = 9'h100 - sizeUDC_io_nextInc;
  assign _T_55 = $unsigned(_T_54);
  assign nextRemainingSlots = _T_55[8:0];
  assign strideDec = io_config_chainRead ? 5'h1 : 5'h10;
  assign _GEN_0 = {{4'd0}, strideDec};
  assign empty = sizeUDC_io_out < _GEN_0;
  assign almostEmpty = sizeUDC_io_nextDec < _GEN_0;
  assign full = remainingSlots < 9'h10;
  assign almostFull = nextRemainingSlots < 9'h10;
  assign _T_64 = ~ full;
  assign writeEn = io_enqVld & _T_64;
  assign _T_65 = ~ empty;
  assign readEn = io_deqVld & _T_65;
  assign _T_101 = readEn & io_config_chainRead;
  assign _T_102 = rptr_io_done_0 ? rptr_io_next_1 : rptr_io_out_1;
  assign nextHeadLocalAddr = io_config_chainRead ? _T_102 : rptr_io_next_1;
  assign _T_154 = readEn ? nextHeadLocalAddr : rptr_io_out_1;
  assign _T_159 = readEn ? rptr_io_next_0 : rptr_io_out_0;
  assign _T_162 = io_config_chainRead ? FF_io_out : 4'h0;
  assign io_deq_0 = MuxN_io_out;
  assign io_deq_1 = mems_0_1_io_rdata;
  assign io_deq_2 = mems_0_2_io_rdata;
  assign io_deq_3 = mems_0_3_io_rdata;
  assign io_deq_4 = mems_0_4_io_rdata;
  assign io_deq_5 = mems_0_5_io_rdata;
  assign io_deq_6 = mems_0_6_io_rdata;
  assign io_deq_7 = mems_0_7_io_rdata;
  assign io_deq_8 = mems_0_8_io_rdata;
  assign io_deq_9 = mems_0_9_io_rdata;
  assign io_deq_10 = mems_0_10_io_rdata;
  assign io_deq_11 = mems_0_11_io_rdata;
  assign io_deq_12 = mems_0_12_io_rdata;
  assign io_deq_13 = mems_0_13_io_rdata;
  assign io_deq_14 = mems_0_14_io_rdata;
  assign io_deq_15 = mems_0_15_io_rdata;
  assign io_full = full;
  assign io_empty = empty;
  assign io_almostFull = almostFull;
  assign io_almostEmpty = almostEmpty;
  assign sizeUDC_io_strideInc = 9'h10;
  assign sizeUDC_io_strideDec = {{4'd0}, strideDec};
  assign sizeUDC_io_inc = writeEn;
  assign sizeUDC_io_dec = readEn;
  assign sizeUDC_clock = clock;
  assign sizeUDC_reset = reset;
  assign wptr_io_enable_0 = 1'h0;
  assign wptr_io_enable_1 = writeEn;
  assign wptr_io_config_chain_0 = 1'h0;
  assign wptr_clock = clock;
  assign wptr_reset = reset;
  assign rptrConfig_chain_0 = io_config_chainRead;
  assign rptr_io_enable_0 = _T_101;
  assign rptr_io_enable_1 = readEn;
  assign rptr_io_config_chain_0 = rptrConfig_chain_0;
  assign rptr_clock = clock;
  assign rptr_reset = reset;
  assign mems_0_0_io_raddr = _T_154[3:0];
  assign mems_0_0_io_wen = writeEn;
  assign mems_0_0_io_waddr = wptr_io_out_1[3:0];
  assign mems_0_0_io_wdata = wdata_0;
  assign mems_0_0_clock = clock;
  assign mems_0_0_reset = reset;
  assign mems_0_1_io_raddr = _T_154[3:0];
  assign mems_0_1_io_wen = writeEn;
  assign mems_0_1_io_waddr = wptr_io_out_1[3:0];
  assign mems_0_1_io_wdata = wdata_1;
  assign mems_0_1_clock = clock;
  assign mems_0_1_reset = reset;
  assign mems_0_2_io_raddr = _T_154[3:0];
  assign mems_0_2_io_wen = writeEn;
  assign mems_0_2_io_waddr = wptr_io_out_1[3:0];
  assign mems_0_2_io_wdata = wdata_2;
  assign mems_0_2_clock = clock;
  assign mems_0_2_reset = reset;
  assign mems_0_3_io_raddr = _T_154[3:0];
  assign mems_0_3_io_wen = writeEn;
  assign mems_0_3_io_waddr = wptr_io_out_1[3:0];
  assign mems_0_3_io_wdata = wdata_3;
  assign mems_0_3_clock = clock;
  assign mems_0_3_reset = reset;
  assign mems_0_4_io_raddr = _T_154[3:0];
  assign mems_0_4_io_wen = writeEn;
  assign mems_0_4_io_waddr = wptr_io_out_1[3:0];
  assign mems_0_4_io_wdata = wdata_4;
  assign mems_0_4_clock = clock;
  assign mems_0_4_reset = reset;
  assign mems_0_5_io_raddr = _T_154[3:0];
  assign mems_0_5_io_wen = writeEn;
  assign mems_0_5_io_waddr = wptr_io_out_1[3:0];
  assign mems_0_5_io_wdata = wdata_5;
  assign mems_0_5_clock = clock;
  assign mems_0_5_reset = reset;
  assign mems_0_6_io_raddr = _T_154[3:0];
  assign mems_0_6_io_wen = writeEn;
  assign mems_0_6_io_waddr = wptr_io_out_1[3:0];
  assign mems_0_6_io_wdata = wdata_6;
  assign mems_0_6_clock = clock;
  assign mems_0_6_reset = reset;
  assign mems_0_7_io_raddr = _T_154[3:0];
  assign mems_0_7_io_wen = writeEn;
  assign mems_0_7_io_waddr = wptr_io_out_1[3:0];
  assign mems_0_7_io_wdata = wdata_7;
  assign mems_0_7_clock = clock;
  assign mems_0_7_reset = reset;
  assign mems_0_8_io_raddr = _T_154[3:0];
  assign mems_0_8_io_wen = writeEn;
  assign mems_0_8_io_waddr = wptr_io_out_1[3:0];
  assign mems_0_8_io_wdata = wdata_8;
  assign mems_0_8_clock = clock;
  assign mems_0_8_reset = reset;
  assign mems_0_9_io_raddr = _T_154[3:0];
  assign mems_0_9_io_wen = writeEn;
  assign mems_0_9_io_waddr = wptr_io_out_1[3:0];
  assign mems_0_9_io_wdata = wdata_9;
  assign mems_0_9_clock = clock;
  assign mems_0_9_reset = reset;
  assign mems_0_10_io_raddr = _T_154[3:0];
  assign mems_0_10_io_wen = writeEn;
  assign mems_0_10_io_waddr = wptr_io_out_1[3:0];
  assign mems_0_10_io_wdata = wdata_10;
  assign mems_0_10_clock = clock;
  assign mems_0_10_reset = reset;
  assign mems_0_11_io_raddr = _T_154[3:0];
  assign mems_0_11_io_wen = writeEn;
  assign mems_0_11_io_waddr = wptr_io_out_1[3:0];
  assign mems_0_11_io_wdata = wdata_11;
  assign mems_0_11_clock = clock;
  assign mems_0_11_reset = reset;
  assign mems_0_12_io_raddr = _T_154[3:0];
  assign mems_0_12_io_wen = writeEn;
  assign mems_0_12_io_waddr = wptr_io_out_1[3:0];
  assign mems_0_12_io_wdata = wdata_12;
  assign mems_0_12_clock = clock;
  assign mems_0_12_reset = reset;
  assign mems_0_13_io_raddr = _T_154[3:0];
  assign mems_0_13_io_wen = writeEn;
  assign mems_0_13_io_waddr = wptr_io_out_1[3:0];
  assign mems_0_13_io_wdata = wdata_13;
  assign mems_0_13_clock = clock;
  assign mems_0_13_reset = reset;
  assign mems_0_14_io_raddr = _T_154[3:0];
  assign mems_0_14_io_wen = writeEn;
  assign mems_0_14_io_waddr = wptr_io_out_1[3:0];
  assign mems_0_14_io_wdata = wdata_14;
  assign mems_0_14_clock = clock;
  assign mems_0_14_reset = reset;
  assign mems_0_15_io_raddr = _T_154[3:0];
  assign mems_0_15_io_wen = writeEn;
  assign mems_0_15_io_waddr = wptr_io_out_1[3:0];
  assign mems_0_15_io_wdata = wdata_15;
  assign mems_0_15_clock = clock;
  assign mems_0_15_reset = reset;
  assign wdata_0 = io_enq_0;
  assign wdata_1 = io_enq_1;
  assign wdata_2 = io_enq_2;
  assign wdata_3 = io_enq_3;
  assign wdata_4 = io_enq_4;
  assign wdata_5 = io_enq_5;
  assign wdata_6 = io_enq_6;
  assign wdata_7 = io_enq_7;
  assign wdata_8 = io_enq_8;
  assign wdata_9 = io_enq_9;
  assign wdata_10 = io_enq_10;
  assign wdata_11 = io_enq_11;
  assign wdata_12 = io_enq_12;
  assign wdata_13 = io_enq_13;
  assign wdata_14 = io_enq_14;
  assign wdata_15 = io_enq_15;
  assign MuxN_io_ins_0 = mems_0_0_io_rdata;
  assign MuxN_io_ins_1 = mems_0_1_io_rdata;
  assign MuxN_io_ins_2 = mems_0_2_io_rdata;
  assign MuxN_io_ins_3 = mems_0_3_io_rdata;
  assign MuxN_io_ins_4 = mems_0_4_io_rdata;
  assign MuxN_io_ins_5 = mems_0_5_io_rdata;
  assign MuxN_io_ins_6 = mems_0_6_io_rdata;
  assign MuxN_io_ins_7 = mems_0_7_io_rdata;
  assign MuxN_io_ins_8 = mems_0_8_io_rdata;
  assign MuxN_io_ins_9 = mems_0_9_io_rdata;
  assign MuxN_io_ins_10 = mems_0_10_io_rdata;
  assign MuxN_io_ins_11 = mems_0_11_io_rdata;
  assign MuxN_io_ins_12 = mems_0_12_io_rdata;
  assign MuxN_io_ins_13 = mems_0_13_io_rdata;
  assign MuxN_io_ins_14 = mems_0_14_io_rdata;
  assign MuxN_io_ins_15 = mems_0_15_io_rdata;
  assign MuxN_io_sel = _T_162;
  assign FF_io_in = _T_159[3:0];
  assign FF_clock = clock;
  assign FF_reset = reset;
endmodule
module SRAM_28(
  input         clock,
  input         reset,
  input  [7:0]  io_raddr,
  input         io_wen,
  input  [7:0]  io_waddr,
  output [15:0] io_rdata
);
  wire [15:0] SRAMVerilogAWS_rdata;
  wire [15:0] SRAMVerilogAWS_wdata;
  wire  SRAMVerilogAWS_flow;
  wire  SRAMVerilogAWS_wen;
  wire  SRAMVerilogAWS_waddrEn;
  wire  SRAMVerilogAWS_raddrEn;
  wire [7:0] SRAMVerilogAWS_waddr;
  wire [7:0] SRAMVerilogAWS_raddr;
  wire  SRAMVerilogAWS_clk;
  wire  _T_8;
  wire  _T_9;
  reg  _T_12;
  reg [31:0] _RAND_0;
  wire [15:0] _T_16;
  wire [15:0] _T_18;
  SRAMVerilogAWS #(.DWIDTH(16), .WORDS(256), .AWIDTH(8)) SRAMVerilogAWS (
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .flow(SRAMVerilogAWS_flow),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_8 = io_raddr == io_waddr;
  assign _T_9 = io_wen & _T_8;
  assign _T_16 = _T_12 ? 16'h0 : SRAMVerilogAWS_rdata;
  assign io_rdata = _T_18;
  assign SRAMVerilogAWS_wdata = 16'h0;
  assign SRAMVerilogAWS_flow = 1'h1;
  assign SRAMVerilogAWS_wen = io_wen;
  assign SRAMVerilogAWS_waddrEn = 1'h1;
  assign SRAMVerilogAWS_raddrEn = 1'h1;
  assign SRAMVerilogAWS_waddr = io_waddr;
  assign SRAMVerilogAWS_raddr = io_raddr;
  assign SRAMVerilogAWS_clk = clock;
  assign _T_18 = _T_16;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_12 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_12 <= 1'h0;
    end else begin
      _T_12 <= _T_9;
    end
  end
endmodule
module MuxN_17(
  input  [15:0] io_ins_0,
  output [15:0] io_out
);
  assign io_out = io_ins_0;
endmodule
module FIFOCore_3(
  input         clock,
  input         reset,
  input         io_enqVld,
  output [15:0] io_deq_0,
  input         io_deqVld,
  input         io_config_chainRead
);
  wire  sizeUDC_clock;
  wire  sizeUDC_reset;
  wire [8:0] sizeUDC_io_strideInc;
  wire [8:0] sizeUDC_io_strideDec;
  wire  sizeUDC_io_inc;
  wire  sizeUDC_io_dec;
  wire [8:0] sizeUDC_io_out;
  wire [8:0] sizeUDC_io_nextInc;
  wire [8:0] sizeUDC_io_nextDec;
  wire [9:0] _T_21;
  wire [9:0] _T_22;
  wire [8:0] remainingSlots;
  wire  empty;
  wire  full;
  wire  _T_34;
  wire  writeEn;
  wire  _T_35;
  wire  readEn;
  wire  wptr_clock;
  wire  wptr_reset;
  wire [8:0] wptr_io_out_0;
  wire [8:0] wptr_io_out_1;
  wire [8:0] wptr_io_next_1;
  wire  wptr_io_enable_0;
  wire  wptr_io_enable_1;
  wire  wptr_io_done_0;
  wire  wptr_io_config_chain_0;
  wire  rptrConfig_chain_0;
  wire  rptr_clock;
  wire  rptr_reset;
  wire [8:0] rptr_io_out_0;
  wire [8:0] rptr_io_out_1;
  wire [8:0] rptr_io_next_1;
  wire  rptr_io_enable_0;
  wire  rptr_io_enable_1;
  wire  rptr_io_done_0;
  wire  rptr_io_config_chain_0;
  wire  _T_71;
  wire [8:0] _T_72;
  wire [8:0] nextHeadLocalAddr;
  wire  mems_0_0_clock;
  wire  mems_0_0_reset;
  wire [7:0] mems_0_0_io_raddr;
  wire  mems_0_0_io_wen;
  wire [7:0] mems_0_0_io_waddr;
  wire [15:0] mems_0_0_io_rdata;
  wire [8:0] _T_79;
  wire [15:0] MuxN_io_ins_0;
  wire [15:0] MuxN_io_out;
  UpDownCtr sizeUDC (
    .clock(sizeUDC_clock),
    .reset(sizeUDC_reset),
    .io_strideInc(sizeUDC_io_strideInc),
    .io_strideDec(sizeUDC_io_strideDec),
    .io_inc(sizeUDC_io_inc),
    .io_dec(sizeUDC_io_dec),
    .io_out(sizeUDC_io_out),
    .io_nextInc(sizeUDC_io_nextInc),
    .io_nextDec(sizeUDC_io_nextDec)
  );
  CounterChainCore wptr (
    .clock(wptr_clock),
    .reset(wptr_reset),
    .io_out_0(wptr_io_out_0),
    .io_out_1(wptr_io_out_1),
    .io_next_1(wptr_io_next_1),
    .io_enable_0(wptr_io_enable_0),
    .io_enable_1(wptr_io_enable_1),
    .io_done_0(wptr_io_done_0),
    .io_config_chain_0(wptr_io_config_chain_0)
  );
  CounterChainCore rptr (
    .clock(rptr_clock),
    .reset(rptr_reset),
    .io_out_0(rptr_io_out_0),
    .io_out_1(rptr_io_out_1),
    .io_next_1(rptr_io_next_1),
    .io_enable_0(rptr_io_enable_0),
    .io_enable_1(rptr_io_enable_1),
    .io_done_0(rptr_io_done_0),
    .io_config_chain_0(rptr_io_config_chain_0)
  );
  SRAM_28 mems_0_0 (
    .clock(mems_0_0_clock),
    .reset(mems_0_0_reset),
    .io_raddr(mems_0_0_io_raddr),
    .io_wen(mems_0_0_io_wen),
    .io_waddr(mems_0_0_io_waddr),
    .io_rdata(mems_0_0_io_rdata)
  );
  MuxN_17 MuxN (
    .io_ins_0(MuxN_io_ins_0),
    .io_out(MuxN_io_out)
  );
  assign _T_21 = 9'h100 - sizeUDC_io_out;
  assign _T_22 = $unsigned(_T_21);
  assign remainingSlots = _T_22[8:0];
  assign empty = sizeUDC_io_out < 9'h1;
  assign full = remainingSlots < 9'h1;
  assign _T_34 = ~ full;
  assign writeEn = io_enqVld & _T_34;
  assign _T_35 = ~ empty;
  assign readEn = io_deqVld & _T_35;
  assign _T_71 = readEn & io_config_chainRead;
  assign _T_72 = rptr_io_done_0 ? rptr_io_next_1 : rptr_io_out_1;
  assign nextHeadLocalAddr = io_config_chainRead ? _T_72 : rptr_io_next_1;
  assign _T_79 = readEn ? nextHeadLocalAddr : rptr_io_out_1;
  assign io_deq_0 = MuxN_io_out;
  assign sizeUDC_io_strideInc = 9'h1;
  assign sizeUDC_io_strideDec = 9'h1;
  assign sizeUDC_io_inc = writeEn;
  assign sizeUDC_io_dec = readEn;
  assign sizeUDC_clock = clock;
  assign sizeUDC_reset = reset;
  assign wptr_io_enable_0 = 1'h0;
  assign wptr_io_enable_1 = writeEn;
  assign wptr_io_config_chain_0 = 1'h0;
  assign wptr_clock = clock;
  assign wptr_reset = reset;
  assign rptrConfig_chain_0 = io_config_chainRead;
  assign rptr_io_enable_0 = _T_71;
  assign rptr_io_enable_1 = readEn;
  assign rptr_io_config_chain_0 = rptrConfig_chain_0;
  assign rptr_clock = clock;
  assign rptr_reset = reset;
  assign mems_0_0_io_raddr = _T_79[7:0];
  assign mems_0_0_io_wen = writeEn;
  assign mems_0_0_io_waddr = wptr_io_out_1[7:0];
  assign mems_0_0_clock = clock;
  assign mems_0_0_reset = reset;
  assign MuxN_io_ins_0 = mems_0_0_io_rdata;
endmodule
module FIFOWidthConvert(
  input         clock,
  input         reset,
  input  [31:0] io_enq_0,
  input  [31:0] io_enq_1,
  input  [31:0] io_enq_2,
  input  [31:0] io_enq_3,
  input  [31:0] io_enq_4,
  input  [31:0] io_enq_5,
  input  [31:0] io_enq_6,
  input  [31:0] io_enq_7,
  input  [31:0] io_enq_8,
  input  [31:0] io_enq_9,
  input  [31:0] io_enq_10,
  input  [31:0] io_enq_11,
  input  [31:0] io_enq_12,
  input  [31:0] io_enq_13,
  input  [31:0] io_enq_14,
  input  [31:0] io_enq_15,
  input         io_enqVld,
  output [31:0] io_deq_0,
  input         io_deqVld,
  output        io_full,
  output        io_empty,
  output        io_almostEmpty,
  output        io_almostFull
);
  wire  FIFOCore_clock;
  wire  FIFOCore_reset;
  wire [31:0] FIFOCore_io_enq_0;
  wire [31:0] FIFOCore_io_enq_1;
  wire [31:0] FIFOCore_io_enq_2;
  wire [31:0] FIFOCore_io_enq_3;
  wire [31:0] FIFOCore_io_enq_4;
  wire [31:0] FIFOCore_io_enq_5;
  wire [31:0] FIFOCore_io_enq_6;
  wire [31:0] FIFOCore_io_enq_7;
  wire [31:0] FIFOCore_io_enq_8;
  wire [31:0] FIFOCore_io_enq_9;
  wire [31:0] FIFOCore_io_enq_10;
  wire [31:0] FIFOCore_io_enq_11;
  wire [31:0] FIFOCore_io_enq_12;
  wire [31:0] FIFOCore_io_enq_13;
  wire [31:0] FIFOCore_io_enq_14;
  wire [31:0] FIFOCore_io_enq_15;
  wire  FIFOCore_io_enqVld;
  wire [31:0] FIFOCore_io_deq_0;
  wire [31:0] FIFOCore_io_deq_1;
  wire [31:0] FIFOCore_io_deq_2;
  wire [31:0] FIFOCore_io_deq_3;
  wire [31:0] FIFOCore_io_deq_4;
  wire [31:0] FIFOCore_io_deq_5;
  wire [31:0] FIFOCore_io_deq_6;
  wire [31:0] FIFOCore_io_deq_7;
  wire [31:0] FIFOCore_io_deq_8;
  wire [31:0] FIFOCore_io_deq_9;
  wire [31:0] FIFOCore_io_deq_10;
  wire [31:0] FIFOCore_io_deq_11;
  wire [31:0] FIFOCore_io_deq_12;
  wire [31:0] FIFOCore_io_deq_13;
  wire [31:0] FIFOCore_io_deq_14;
  wire [31:0] FIFOCore_io_deq_15;
  wire  FIFOCore_io_deqVld;
  wire  FIFOCore_io_full;
  wire  FIFOCore_io_empty;
  wire  FIFOCore_io_almostFull;
  wire  FIFOCore_io_almostEmpty;
  wire  FIFOCore_io_config_chainRead;
  wire  FIFOCore_1_clock;
  wire  FIFOCore_1_reset;
  wire  FIFOCore_1_io_enqVld;
  wire [15:0] FIFOCore_1_io_deq_0;
  wire  FIFOCore_1_io_deqVld;
  wire  FIFOCore_1_io_config_chainRead;
  wire [63:0] _T_42;
  wire [95:0] _T_43;
  wire [127:0] _T_44;
  wire [159:0] _T_45;
  wire [191:0] _T_46;
  wire [223:0] _T_47;
  wire [255:0] _T_48;
  wire [287:0] _T_49;
  wire [319:0] _T_50;
  wire [351:0] _T_51;
  wire [383:0] _T_52;
  wire [415:0] _T_53;
  wire [447:0] _T_54;
  wire [479:0] _T_55;
  wire [511:0] _T_56;
  wire [31:0] _T_57;
  wire [31:0] _T_58;
  wire [31:0] _T_59;
  wire [31:0] _T_60;
  wire [31:0] _T_61;
  wire [31:0] _T_62;
  wire [31:0] _T_63;
  wire [31:0] _T_64;
  wire [31:0] _T_65;
  wire [31:0] _T_66;
  wire [31:0] _T_67;
  wire [31:0] _T_68;
  wire [31:0] _T_69;
  wire [31:0] _T_70;
  wire [31:0] _T_71;
  wire [31:0] _T_72;
  wire [31:0] _T_75_0;
  wire [31:0] _T_75_1;
  wire [31:0] _T_75_2;
  wire [31:0] _T_75_3;
  wire [31:0] _T_75_4;
  wire [31:0] _T_75_5;
  wire [31:0] _T_75_6;
  wire [31:0] _T_75_7;
  wire [31:0] _T_75_8;
  wire [31:0] _T_75_9;
  wire [31:0] _T_75_10;
  wire [31:0] _T_75_11;
  wire [31:0] _T_75_12;
  wire [31:0] _T_75_13;
  wire [31:0] _T_75_14;
  wire [31:0] _T_75_15;
  wire [31:0] _T_96_0;
  wire [31:0] _T_103_0;
  FIFOCore_2 FIFOCore (
    .clock(FIFOCore_clock),
    .reset(FIFOCore_reset),
    .io_enq_0(FIFOCore_io_enq_0),
    .io_enq_1(FIFOCore_io_enq_1),
    .io_enq_2(FIFOCore_io_enq_2),
    .io_enq_3(FIFOCore_io_enq_3),
    .io_enq_4(FIFOCore_io_enq_4),
    .io_enq_5(FIFOCore_io_enq_5),
    .io_enq_6(FIFOCore_io_enq_6),
    .io_enq_7(FIFOCore_io_enq_7),
    .io_enq_8(FIFOCore_io_enq_8),
    .io_enq_9(FIFOCore_io_enq_9),
    .io_enq_10(FIFOCore_io_enq_10),
    .io_enq_11(FIFOCore_io_enq_11),
    .io_enq_12(FIFOCore_io_enq_12),
    .io_enq_13(FIFOCore_io_enq_13),
    .io_enq_14(FIFOCore_io_enq_14),
    .io_enq_15(FIFOCore_io_enq_15),
    .io_enqVld(FIFOCore_io_enqVld),
    .io_deq_0(FIFOCore_io_deq_0),
    .io_deq_1(FIFOCore_io_deq_1),
    .io_deq_2(FIFOCore_io_deq_2),
    .io_deq_3(FIFOCore_io_deq_3),
    .io_deq_4(FIFOCore_io_deq_4),
    .io_deq_5(FIFOCore_io_deq_5),
    .io_deq_6(FIFOCore_io_deq_6),
    .io_deq_7(FIFOCore_io_deq_7),
    .io_deq_8(FIFOCore_io_deq_8),
    .io_deq_9(FIFOCore_io_deq_9),
    .io_deq_10(FIFOCore_io_deq_10),
    .io_deq_11(FIFOCore_io_deq_11),
    .io_deq_12(FIFOCore_io_deq_12),
    .io_deq_13(FIFOCore_io_deq_13),
    .io_deq_14(FIFOCore_io_deq_14),
    .io_deq_15(FIFOCore_io_deq_15),
    .io_deqVld(FIFOCore_io_deqVld),
    .io_full(FIFOCore_io_full),
    .io_empty(FIFOCore_io_empty),
    .io_almostFull(FIFOCore_io_almostFull),
    .io_almostEmpty(FIFOCore_io_almostEmpty),
    .io_config_chainRead(FIFOCore_io_config_chainRead)
  );
  FIFOCore_3 FIFOCore_1 (
    .clock(FIFOCore_1_clock),
    .reset(FIFOCore_1_reset),
    .io_enqVld(FIFOCore_1_io_enqVld),
    .io_deq_0(FIFOCore_1_io_deq_0),
    .io_deqVld(FIFOCore_1_io_deqVld),
    .io_config_chainRead(FIFOCore_1_io_config_chainRead)
  );
  assign _T_42 = {io_enq_15,io_enq_14};
  assign _T_43 = {_T_42,io_enq_13};
  assign _T_44 = {_T_43,io_enq_12};
  assign _T_45 = {_T_44,io_enq_11};
  assign _T_46 = {_T_45,io_enq_10};
  assign _T_47 = {_T_46,io_enq_9};
  assign _T_48 = {_T_47,io_enq_8};
  assign _T_49 = {_T_48,io_enq_7};
  assign _T_50 = {_T_49,io_enq_6};
  assign _T_51 = {_T_50,io_enq_5};
  assign _T_52 = {_T_51,io_enq_4};
  assign _T_53 = {_T_52,io_enq_3};
  assign _T_54 = {_T_53,io_enq_2};
  assign _T_55 = {_T_54,io_enq_1};
  assign _T_56 = {_T_55,io_enq_0};
  assign _T_57 = _T_56[31:0];
  assign _T_58 = _T_56[63:32];
  assign _T_59 = _T_56[95:64];
  assign _T_60 = _T_56[127:96];
  assign _T_61 = _T_56[159:128];
  assign _T_62 = _T_56[191:160];
  assign _T_63 = _T_56[223:192];
  assign _T_64 = _T_56[255:224];
  assign _T_65 = _T_56[287:256];
  assign _T_66 = _T_56[319:288];
  assign _T_67 = _T_56[351:320];
  assign _T_68 = _T_56[383:352];
  assign _T_69 = _T_56[415:384];
  assign _T_70 = _T_56[447:416];
  assign _T_71 = _T_56[479:448];
  assign _T_72 = _T_56[511:480];
  assign io_deq_0 = _T_103_0;
  assign io_full = FIFOCore_io_full;
  assign io_empty = FIFOCore_io_empty;
  assign io_almostEmpty = FIFOCore_io_almostEmpty;
  assign io_almostFull = FIFOCore_io_almostFull;
  assign FIFOCore_io_enq_0 = _T_75_0;
  assign FIFOCore_io_enq_1 = _T_75_1;
  assign FIFOCore_io_enq_2 = _T_75_2;
  assign FIFOCore_io_enq_3 = _T_75_3;
  assign FIFOCore_io_enq_4 = _T_75_4;
  assign FIFOCore_io_enq_5 = _T_75_5;
  assign FIFOCore_io_enq_6 = _T_75_6;
  assign FIFOCore_io_enq_7 = _T_75_7;
  assign FIFOCore_io_enq_8 = _T_75_8;
  assign FIFOCore_io_enq_9 = _T_75_9;
  assign FIFOCore_io_enq_10 = _T_75_10;
  assign FIFOCore_io_enq_11 = _T_75_11;
  assign FIFOCore_io_enq_12 = _T_75_12;
  assign FIFOCore_io_enq_13 = _T_75_13;
  assign FIFOCore_io_enq_14 = _T_75_14;
  assign FIFOCore_io_enq_15 = _T_75_15;
  assign FIFOCore_io_enqVld = io_enqVld;
  assign FIFOCore_io_deqVld = io_deqVld;
  assign FIFOCore_io_config_chainRead = 1'h1;
  assign FIFOCore_clock = clock;
  assign FIFOCore_reset = reset;
  assign FIFOCore_1_io_enqVld = io_enqVld;
  assign FIFOCore_1_io_deqVld = 1'h0;
  assign FIFOCore_1_io_config_chainRead = 1'h1;
  assign FIFOCore_1_clock = clock;
  assign FIFOCore_1_reset = reset;
  assign _T_75_0 = _T_57;
  assign _T_75_1 = _T_58;
  assign _T_75_2 = _T_59;
  assign _T_75_3 = _T_60;
  assign _T_75_4 = _T_61;
  assign _T_75_5 = _T_62;
  assign _T_75_6 = _T_63;
  assign _T_75_7 = _T_64;
  assign _T_75_8 = _T_65;
  assign _T_75_9 = _T_66;
  assign _T_75_10 = _T_67;
  assign _T_75_11 = _T_68;
  assign _T_75_12 = _T_69;
  assign _T_75_13 = _T_70;
  assign _T_75_14 = _T_71;
  assign _T_75_15 = _T_72;
  assign _T_96_0 = FIFOCore_io_deq_0;
  assign _T_103_0 = _T_96_0;
endmodule
module RetimeWrapper_622(
  input          clock,
  input          reset,
  input  [511:0] io_in,
  output [511:0] io_out
);
  wire [511:0] sr_out;
  wire [511:0] sr_in;
  wire  sr_flow;
  wire  sr_reset;
  wire  sr_clock;
  RetimeShiftRegister #(.WIDTH(512), .STAGES(1)) sr (
    .out(sr_out),
    .in(sr_in),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out;
  assign sr_in = io_in;
  assign sr_flow = 1'h1;
  assign sr_reset = reset;
  assign sr_clock = clock;
endmodule
module FF_180(
  input          clock,
  input          reset,
  input  [511:0] io_in,
  output [511:0] io_out,
  input          io_enable
);
  wire [511:0] d;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire [511:0] RetimeWrapper_io_in;
  wire [511:0] RetimeWrapper_io_out;
  wire [511:0] _T_11;
  wire [511:0] _GEN_1;
  RetimeWrapper_622 RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _GEN_1 = io_enable ? io_in : _T_11;
  assign io_out = _T_11;
  assign d = _GEN_1;
  assign RetimeWrapper_io_in = d;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_11 = RetimeWrapper_io_out;
endmodule
module FIFOWidthConvert_1(
  input         clock,
  input         reset,
  input         io_enqVld,
  output [31:0] io_deq_0,
  output [31:0] io_deq_1,
  output [31:0] io_deq_2,
  output [31:0] io_deq_3,
  output [31:0] io_deq_4,
  output [31:0] io_deq_5,
  output [31:0] io_deq_6,
  output [31:0] io_deq_7,
  output [31:0] io_deq_8,
  output [31:0] io_deq_9,
  output [31:0] io_deq_10,
  output [31:0] io_deq_11,
  output [31:0] io_deq_12,
  output [31:0] io_deq_13,
  output [31:0] io_deq_14,
  output [31:0] io_deq_15,
  output [63:0] io_deqStrb,
  input         io_deqVld,
  output        io_full,
  output        io_empty,
  output        io_almostEmpty,
  output        io_almostFull
);
  wire  FIFOCore_clock;
  wire  FIFOCore_reset;
  wire [31:0] FIFOCore_io_enq_0;
  wire [31:0] FIFOCore_io_enq_1;
  wire [31:0] FIFOCore_io_enq_2;
  wire [31:0] FIFOCore_io_enq_3;
  wire [31:0] FIFOCore_io_enq_4;
  wire [31:0] FIFOCore_io_enq_5;
  wire [31:0] FIFOCore_io_enq_6;
  wire [31:0] FIFOCore_io_enq_7;
  wire [31:0] FIFOCore_io_enq_8;
  wire [31:0] FIFOCore_io_enq_9;
  wire [31:0] FIFOCore_io_enq_10;
  wire [31:0] FIFOCore_io_enq_11;
  wire [31:0] FIFOCore_io_enq_12;
  wire [31:0] FIFOCore_io_enq_13;
  wire [31:0] FIFOCore_io_enq_14;
  wire [31:0] FIFOCore_io_enq_15;
  wire  FIFOCore_io_enqVld;
  wire [31:0] FIFOCore_io_deq_0;
  wire [31:0] FIFOCore_io_deq_1;
  wire [31:0] FIFOCore_io_deq_2;
  wire [31:0] FIFOCore_io_deq_3;
  wire [31:0] FIFOCore_io_deq_4;
  wire [31:0] FIFOCore_io_deq_5;
  wire [31:0] FIFOCore_io_deq_6;
  wire [31:0] FIFOCore_io_deq_7;
  wire [31:0] FIFOCore_io_deq_8;
  wire [31:0] FIFOCore_io_deq_9;
  wire [31:0] FIFOCore_io_deq_10;
  wire [31:0] FIFOCore_io_deq_11;
  wire [31:0] FIFOCore_io_deq_12;
  wire [31:0] FIFOCore_io_deq_13;
  wire [31:0] FIFOCore_io_deq_14;
  wire [31:0] FIFOCore_io_deq_15;
  wire  FIFOCore_io_deqVld;
  wire  FIFOCore_io_full;
  wire  FIFOCore_io_empty;
  wire  FIFOCore_io_almostFull;
  wire  FIFOCore_io_almostEmpty;
  wire  FIFOCore_io_config_chainRead;
  wire  FIFOCore_1_clock;
  wire  FIFOCore_1_reset;
  wire  FIFOCore_1_io_enqVld;
  wire [15:0] FIFOCore_1_io_deq_0;
  wire  FIFOCore_1_io_deqVld;
  wire  FIFOCore_1_io_config_chainRead;
  wire  _T_57;
  wire  _T_61;
  wire  _T_65;
  wire  _T_69;
  wire  _T_73;
  wire  _T_77;
  wire  _T_81;
  wire  _T_85;
  wire  _T_89;
  wire  _T_93;
  wire  _T_97;
  wire  _T_101;
  wire  _T_105;
  wire  _T_109;
  wire  _T_113;
  wire  _T_117;
  wire  _T_123_0;
  wire  _T_123_1;
  wire  _T_123_2;
  wire  _T_123_3;
  wire  _T_123_4;
  wire  _T_123_5;
  wire  _T_123_6;
  wire  _T_123_7;
  wire  _T_123_8;
  wire  _T_123_9;
  wire  _T_123_10;
  wire  _T_123_11;
  wire  _T_123_12;
  wire  _T_123_13;
  wire  _T_123_14;
  wire  _T_123_15;
  wire  _T_123_16;
  wire  _T_123_17;
  wire  _T_123_18;
  wire  _T_123_19;
  wire  _T_123_20;
  wire  _T_123_21;
  wire  _T_123_22;
  wire  _T_123_23;
  wire  _T_123_24;
  wire  _T_123_25;
  wire  _T_123_26;
  wire  _T_123_27;
  wire  _T_123_28;
  wire  _T_123_29;
  wire  _T_123_30;
  wire  _T_123_31;
  wire  _T_123_32;
  wire  _T_123_33;
  wire  _T_123_34;
  wire  _T_123_35;
  wire  _T_123_36;
  wire  _T_123_37;
  wire  _T_123_38;
  wire  _T_123_39;
  wire  _T_123_40;
  wire  _T_123_41;
  wire  _T_123_42;
  wire  _T_123_43;
  wire  _T_123_44;
  wire  _T_123_45;
  wire  _T_123_46;
  wire  _T_123_47;
  wire  _T_123_48;
  wire  _T_123_49;
  wire  _T_123_50;
  wire  _T_123_51;
  wire  _T_123_52;
  wire  _T_123_53;
  wire  _T_123_54;
  wire  _T_123_55;
  wire  _T_123_56;
  wire  _T_123_57;
  wire  _T_123_58;
  wire  _T_123_59;
  wire  _T_123_60;
  wire  _T_123_61;
  wire  _T_123_62;
  wire  _T_123_63;
  wire [1:0] _T_190;
  wire [2:0] _T_191;
  wire [3:0] _T_192;
  wire [4:0] _T_193;
  wire [5:0] _T_194;
  wire [6:0] _T_195;
  wire [7:0] _T_196;
  wire [8:0] _T_197;
  wire [9:0] _T_198;
  wire [10:0] _T_199;
  wire [11:0] _T_200;
  wire [12:0] _T_201;
  wire [13:0] _T_202;
  wire [14:0] _T_203;
  wire [15:0] _T_204;
  wire [16:0] _T_205;
  wire [17:0] _T_206;
  wire [18:0] _T_207;
  wire [19:0] _T_208;
  wire [20:0] _T_209;
  wire [21:0] _T_210;
  wire [22:0] _T_211;
  wire [23:0] _T_212;
  wire [24:0] _T_213;
  wire [25:0] _T_214;
  wire [26:0] _T_215;
  wire [27:0] _T_216;
  wire [28:0] _T_217;
  wire [29:0] _T_218;
  wire [30:0] _T_219;
  wire [31:0] _T_220;
  wire [32:0] _T_221;
  wire [33:0] _T_222;
  wire [34:0] _T_223;
  wire [35:0] _T_224;
  wire [36:0] _T_225;
  wire [37:0] _T_226;
  wire [38:0] _T_227;
  wire [39:0] _T_228;
  wire [40:0] _T_229;
  wire [41:0] _T_230;
  wire [42:0] _T_231;
  wire [43:0] _T_232;
  wire [44:0] _T_233;
  wire [45:0] _T_234;
  wire [46:0] _T_235;
  wire [47:0] _T_236;
  wire [48:0] _T_237;
  wire [49:0] _T_238;
  wire [50:0] _T_239;
  wire [51:0] _T_240;
  wire [52:0] _T_241;
  wire [53:0] _T_242;
  wire [54:0] _T_243;
  wire [55:0] _T_244;
  wire [56:0] _T_245;
  wire [57:0] _T_246;
  wire [58:0] _T_247;
  wire [59:0] _T_248;
  wire [60:0] _T_249;
  wire [61:0] _T_250;
  wire [62:0] _T_251;
  wire [63:0] _T_252;
  FIFOCore_2 FIFOCore (
    .clock(FIFOCore_clock),
    .reset(FIFOCore_reset),
    .io_enq_0(FIFOCore_io_enq_0),
    .io_enq_1(FIFOCore_io_enq_1),
    .io_enq_2(FIFOCore_io_enq_2),
    .io_enq_3(FIFOCore_io_enq_3),
    .io_enq_4(FIFOCore_io_enq_4),
    .io_enq_5(FIFOCore_io_enq_5),
    .io_enq_6(FIFOCore_io_enq_6),
    .io_enq_7(FIFOCore_io_enq_7),
    .io_enq_8(FIFOCore_io_enq_8),
    .io_enq_9(FIFOCore_io_enq_9),
    .io_enq_10(FIFOCore_io_enq_10),
    .io_enq_11(FIFOCore_io_enq_11),
    .io_enq_12(FIFOCore_io_enq_12),
    .io_enq_13(FIFOCore_io_enq_13),
    .io_enq_14(FIFOCore_io_enq_14),
    .io_enq_15(FIFOCore_io_enq_15),
    .io_enqVld(FIFOCore_io_enqVld),
    .io_deq_0(FIFOCore_io_deq_0),
    .io_deq_1(FIFOCore_io_deq_1),
    .io_deq_2(FIFOCore_io_deq_2),
    .io_deq_3(FIFOCore_io_deq_3),
    .io_deq_4(FIFOCore_io_deq_4),
    .io_deq_5(FIFOCore_io_deq_5),
    .io_deq_6(FIFOCore_io_deq_6),
    .io_deq_7(FIFOCore_io_deq_7),
    .io_deq_8(FIFOCore_io_deq_8),
    .io_deq_9(FIFOCore_io_deq_9),
    .io_deq_10(FIFOCore_io_deq_10),
    .io_deq_11(FIFOCore_io_deq_11),
    .io_deq_12(FIFOCore_io_deq_12),
    .io_deq_13(FIFOCore_io_deq_13),
    .io_deq_14(FIFOCore_io_deq_14),
    .io_deq_15(FIFOCore_io_deq_15),
    .io_deqVld(FIFOCore_io_deqVld),
    .io_full(FIFOCore_io_full),
    .io_empty(FIFOCore_io_empty),
    .io_almostFull(FIFOCore_io_almostFull),
    .io_almostEmpty(FIFOCore_io_almostEmpty),
    .io_config_chainRead(FIFOCore_io_config_chainRead)
  );
  FIFOCore_3 FIFOCore_1 (
    .clock(FIFOCore_1_clock),
    .reset(FIFOCore_1_reset),
    .io_enqVld(FIFOCore_1_io_enqVld),
    .io_deq_0(FIFOCore_1_io_deq_0),
    .io_deqVld(FIFOCore_1_io_deqVld),
    .io_config_chainRead(FIFOCore_1_io_config_chainRead)
  );
  assign _T_57 = FIFOCore_1_io_deq_0[0];
  assign _T_61 = FIFOCore_1_io_deq_0[1];
  assign _T_65 = FIFOCore_1_io_deq_0[2];
  assign _T_69 = FIFOCore_1_io_deq_0[3];
  assign _T_73 = FIFOCore_1_io_deq_0[4];
  assign _T_77 = FIFOCore_1_io_deq_0[5];
  assign _T_81 = FIFOCore_1_io_deq_0[6];
  assign _T_85 = FIFOCore_1_io_deq_0[7];
  assign _T_89 = FIFOCore_1_io_deq_0[8];
  assign _T_93 = FIFOCore_1_io_deq_0[9];
  assign _T_97 = FIFOCore_1_io_deq_0[10];
  assign _T_101 = FIFOCore_1_io_deq_0[11];
  assign _T_105 = FIFOCore_1_io_deq_0[12];
  assign _T_109 = FIFOCore_1_io_deq_0[13];
  assign _T_113 = FIFOCore_1_io_deq_0[14];
  assign _T_117 = FIFOCore_1_io_deq_0[15];
  assign _T_190 = {_T_123_0,_T_123_1};
  assign _T_191 = {_T_190,_T_123_2};
  assign _T_192 = {_T_191,_T_123_3};
  assign _T_193 = {_T_192,_T_123_4};
  assign _T_194 = {_T_193,_T_123_5};
  assign _T_195 = {_T_194,_T_123_6};
  assign _T_196 = {_T_195,_T_123_7};
  assign _T_197 = {_T_196,_T_123_8};
  assign _T_198 = {_T_197,_T_123_9};
  assign _T_199 = {_T_198,_T_123_10};
  assign _T_200 = {_T_199,_T_123_11};
  assign _T_201 = {_T_200,_T_123_12};
  assign _T_202 = {_T_201,_T_123_13};
  assign _T_203 = {_T_202,_T_123_14};
  assign _T_204 = {_T_203,_T_123_15};
  assign _T_205 = {_T_204,_T_123_16};
  assign _T_206 = {_T_205,_T_123_17};
  assign _T_207 = {_T_206,_T_123_18};
  assign _T_208 = {_T_207,_T_123_19};
  assign _T_209 = {_T_208,_T_123_20};
  assign _T_210 = {_T_209,_T_123_21};
  assign _T_211 = {_T_210,_T_123_22};
  assign _T_212 = {_T_211,_T_123_23};
  assign _T_213 = {_T_212,_T_123_24};
  assign _T_214 = {_T_213,_T_123_25};
  assign _T_215 = {_T_214,_T_123_26};
  assign _T_216 = {_T_215,_T_123_27};
  assign _T_217 = {_T_216,_T_123_28};
  assign _T_218 = {_T_217,_T_123_29};
  assign _T_219 = {_T_218,_T_123_30};
  assign _T_220 = {_T_219,_T_123_31};
  assign _T_221 = {_T_220,_T_123_32};
  assign _T_222 = {_T_221,_T_123_33};
  assign _T_223 = {_T_222,_T_123_34};
  assign _T_224 = {_T_223,_T_123_35};
  assign _T_225 = {_T_224,_T_123_36};
  assign _T_226 = {_T_225,_T_123_37};
  assign _T_227 = {_T_226,_T_123_38};
  assign _T_228 = {_T_227,_T_123_39};
  assign _T_229 = {_T_228,_T_123_40};
  assign _T_230 = {_T_229,_T_123_41};
  assign _T_231 = {_T_230,_T_123_42};
  assign _T_232 = {_T_231,_T_123_43};
  assign _T_233 = {_T_232,_T_123_44};
  assign _T_234 = {_T_233,_T_123_45};
  assign _T_235 = {_T_234,_T_123_46};
  assign _T_236 = {_T_235,_T_123_47};
  assign _T_237 = {_T_236,_T_123_48};
  assign _T_238 = {_T_237,_T_123_49};
  assign _T_239 = {_T_238,_T_123_50};
  assign _T_240 = {_T_239,_T_123_51};
  assign _T_241 = {_T_240,_T_123_52};
  assign _T_242 = {_T_241,_T_123_53};
  assign _T_243 = {_T_242,_T_123_54};
  assign _T_244 = {_T_243,_T_123_55};
  assign _T_245 = {_T_244,_T_123_56};
  assign _T_246 = {_T_245,_T_123_57};
  assign _T_247 = {_T_246,_T_123_58};
  assign _T_248 = {_T_247,_T_123_59};
  assign _T_249 = {_T_248,_T_123_60};
  assign _T_250 = {_T_249,_T_123_61};
  assign _T_251 = {_T_250,_T_123_62};
  assign _T_252 = {_T_251,_T_123_63};
  assign io_deq_0 = FIFOCore_io_deq_0;
  assign io_deq_1 = FIFOCore_io_deq_1;
  assign io_deq_2 = FIFOCore_io_deq_2;
  assign io_deq_3 = FIFOCore_io_deq_3;
  assign io_deq_4 = FIFOCore_io_deq_4;
  assign io_deq_5 = FIFOCore_io_deq_5;
  assign io_deq_6 = FIFOCore_io_deq_6;
  assign io_deq_7 = FIFOCore_io_deq_7;
  assign io_deq_8 = FIFOCore_io_deq_8;
  assign io_deq_9 = FIFOCore_io_deq_9;
  assign io_deq_10 = FIFOCore_io_deq_10;
  assign io_deq_11 = FIFOCore_io_deq_11;
  assign io_deq_12 = FIFOCore_io_deq_12;
  assign io_deq_13 = FIFOCore_io_deq_13;
  assign io_deq_14 = FIFOCore_io_deq_14;
  assign io_deq_15 = FIFOCore_io_deq_15;
  assign io_deqStrb = _T_252;
  assign io_full = FIFOCore_io_full;
  assign io_empty = FIFOCore_io_empty;
  assign io_almostEmpty = FIFOCore_io_almostEmpty;
  assign io_almostFull = FIFOCore_io_almostFull;
  assign FIFOCore_io_enq_0 = 32'h0;
  assign FIFOCore_io_enq_1 = 32'h0;
  assign FIFOCore_io_enq_2 = 32'h0;
  assign FIFOCore_io_enq_3 = 32'h0;
  assign FIFOCore_io_enq_4 = 32'h0;
  assign FIFOCore_io_enq_5 = 32'h0;
  assign FIFOCore_io_enq_6 = 32'h0;
  assign FIFOCore_io_enq_7 = 32'h0;
  assign FIFOCore_io_enq_8 = 32'h0;
  assign FIFOCore_io_enq_9 = 32'h0;
  assign FIFOCore_io_enq_10 = 32'h0;
  assign FIFOCore_io_enq_11 = 32'h0;
  assign FIFOCore_io_enq_12 = 32'h0;
  assign FIFOCore_io_enq_13 = 32'h0;
  assign FIFOCore_io_enq_14 = 32'h0;
  assign FIFOCore_io_enq_15 = 32'h0;
  assign FIFOCore_io_enqVld = 1'h0;
  assign FIFOCore_io_deqVld = io_deqVld;
  assign FIFOCore_io_config_chainRead = 1'h0;
  assign FIFOCore_clock = clock;
  assign FIFOCore_reset = reset;
  assign FIFOCore_1_io_enqVld = 1'h0;
  assign FIFOCore_1_io_deqVld = io_deqVld;
  assign FIFOCore_1_io_config_chainRead = 1'h0;
  assign FIFOCore_1_clock = clock;
  assign FIFOCore_1_reset = reset;
  assign _T_123_0 = _T_117;
  assign _T_123_1 = _T_117;
  assign _T_123_2 = _T_117;
  assign _T_123_3 = _T_117;
  assign _T_123_4 = _T_113;
  assign _T_123_5 = _T_113;
  assign _T_123_6 = _T_113;
  assign _T_123_7 = _T_113;
  assign _T_123_8 = _T_109;
  assign _T_123_9 = _T_109;
  assign _T_123_10 = _T_109;
  assign _T_123_11 = _T_109;
  assign _T_123_12 = _T_105;
  assign _T_123_13 = _T_105;
  assign _T_123_14 = _T_105;
  assign _T_123_15 = _T_105;
  assign _T_123_16 = _T_101;
  assign _T_123_17 = _T_101;
  assign _T_123_18 = _T_101;
  assign _T_123_19 = _T_101;
  assign _T_123_20 = _T_97;
  assign _T_123_21 = _T_97;
  assign _T_123_22 = _T_97;
  assign _T_123_23 = _T_97;
  assign _T_123_24 = _T_93;
  assign _T_123_25 = _T_93;
  assign _T_123_26 = _T_93;
  assign _T_123_27 = _T_93;
  assign _T_123_28 = _T_89;
  assign _T_123_29 = _T_89;
  assign _T_123_30 = _T_89;
  assign _T_123_31 = _T_89;
  assign _T_123_32 = _T_85;
  assign _T_123_33 = _T_85;
  assign _T_123_34 = _T_85;
  assign _T_123_35 = _T_85;
  assign _T_123_36 = _T_81;
  assign _T_123_37 = _T_81;
  assign _T_123_38 = _T_81;
  assign _T_123_39 = _T_81;
  assign _T_123_40 = _T_77;
  assign _T_123_41 = _T_77;
  assign _T_123_42 = _T_77;
  assign _T_123_43 = _T_77;
  assign _T_123_44 = _T_73;
  assign _T_123_45 = _T_73;
  assign _T_123_46 = _T_73;
  assign _T_123_47 = _T_73;
  assign _T_123_48 = _T_69;
  assign _T_123_49 = _T_69;
  assign _T_123_50 = _T_69;
  assign _T_123_51 = _T_69;
  assign _T_123_52 = _T_65;
  assign _T_123_53 = _T_65;
  assign _T_123_54 = _T_65;
  assign _T_123_55 = _T_65;
  assign _T_123_56 = _T_61;
  assign _T_123_57 = _T_61;
  assign _T_123_58 = _T_61;
  assign _T_123_59 = _T_61;
  assign _T_123_60 = _T_57;
  assign _T_123_61 = _T_57;
  assign _T_123_62 = _T_57;
  assign _T_123_63 = _T_57;
endmodule
module FIFOCounter(
  input   clock,
  input   reset,
  input   io_enqVld,
  output  io_full,
  output  io_empty
);
  wire  sizeUDC_clock;
  wire  sizeUDC_reset;
  wire [8:0] sizeUDC_io_strideInc;
  wire [8:0] sizeUDC_io_strideDec;
  wire  sizeUDC_io_inc;
  wire  sizeUDC_io_dec;
  wire [8:0] sizeUDC_io_out;
  wire [8:0] sizeUDC_io_nextInc;
  wire [8:0] sizeUDC_io_nextDec;
  wire [9:0] _T_21;
  wire [9:0] _T_22;
  wire [8:0] remainingSlots;
  wire  empty;
  wire  full;
  wire  _T_34;
  wire  writeEn;
  UpDownCtr sizeUDC (
    .clock(sizeUDC_clock),
    .reset(sizeUDC_reset),
    .io_strideInc(sizeUDC_io_strideInc),
    .io_strideDec(sizeUDC_io_strideDec),
    .io_inc(sizeUDC_io_inc),
    .io_dec(sizeUDC_io_dec),
    .io_out(sizeUDC_io_out),
    .io_nextInc(sizeUDC_io_nextInc),
    .io_nextDec(sizeUDC_io_nextDec)
  );
  assign _T_21 = 9'h100 - sizeUDC_io_out;
  assign _T_22 = $unsigned(_T_21);
  assign remainingSlots = _T_22[8:0];
  assign empty = sizeUDC_io_out < 9'h1;
  assign full = remainingSlots < 9'h1;
  assign _T_34 = ~ full;
  assign writeEn = io_enqVld & _T_34;
  assign io_full = full;
  assign io_empty = empty;
  assign sizeUDC_io_strideInc = 9'h1;
  assign sizeUDC_io_strideDec = 9'h1;
  assign sizeUDC_io_inc = writeEn;
  assign sizeUDC_io_dec = 1'h0;
  assign sizeUDC_clock = clock;
  assign sizeUDC_reset = reset;
endmodule
module RetimeWrapper_706(
  input        clock,
  input        reset,
  input  [7:0] io_in,
  output [7:0] io_out
);
  wire [7:0] sr_out;
  wire [7:0] sr_in;
  wire  sr_flow;
  wire  sr_reset;
  wire  sr_clock;
  RetimeShiftRegister #(.WIDTH(8), .STAGES(1)) sr (
    .out(sr_out),
    .in(sr_in),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out;
  assign sr_in = io_in;
  assign sr_flow = 1'h1;
  assign sr_reset = reset;
  assign sr_clock = clock;
endmodule
module FF_265(
  input        clock,
  input        reset,
  input  [7:0] io_in,
  output [7:0] io_out,
  input        io_enable
);
  wire [7:0] d;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire [7:0] RetimeWrapper_io_in;
  wire [7:0] RetimeWrapper_io_out;
  wire [7:0] _T_11;
  wire [7:0] _GEN_1;
  RetimeWrapper_706 RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _GEN_1 = io_enable ? io_in : _T_11;
  assign io_out = _T_11;
  assign d = _GEN_1;
  assign RetimeWrapper_io_in = d;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_11 = RetimeWrapper_io_out;
endmodule
module FF_266(
  input        clock,
  input        reset,
  input  [2:0] io_in,
  output [2:0] io_out,
  input        io_enable
);
  wire [2:0] d;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire [2:0] RetimeWrapper_io_in;
  wire [2:0] RetimeWrapper_io_out;
  wire [2:0] _T_11;
  wire [2:0] _GEN_1;
  RetimeWrapper_106 RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _GEN_1 = io_enable ? io_in : _T_11;
  assign io_out = _T_11;
  assign d = _GEN_1;
  assign RetimeWrapper_io_in = d;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_11 = RetimeWrapper_io_out;
endmodule
module FF_268(
  input        clock,
  input        reset,
  input  [1:0] io_in,
  output [1:0] io_out,
  input        io_enable
);
  wire [1:0] d;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire [1:0] RetimeWrapper_io_in;
  wire [1:0] RetimeWrapper_io_out;
  wire [1:0] _T_11;
  wire [1:0] _GEN_1;
  RetimeWrapper_182 RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _GEN_1 = io_enable ? io_in : _T_11;
  assign io_out = _T_11;
  assign d = _GEN_1;
  assign RetimeWrapper_io_in = d;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_11 = RetimeWrapper_io_out;
endmodule
module MAGCore(
  input          clock,
  input          reset,
  input          io_enable,
  input          io_reset,
  output         io_app_loads_0_cmd_ready,
  input          io_app_loads_0_cmd_valid,
  input  [63:0]  io_app_loads_0_cmd_bits_addr,
  input          io_app_loads_0_cmd_bits_isWr,
  input  [15:0]  io_app_loads_0_cmd_bits_size,
  input          io_app_loads_0_rdata_ready,
  output         io_app_loads_0_rdata_valid,
  output [31:0]  io_app_loads_0_rdata_bits_0,
  input          io_dram_cmd_ready,
  output         io_dram_cmd_valid,
  output [63:0]  io_dram_cmd_bits_addr,
  output [31:0]  io_dram_cmd_bits_size,
  output         io_dram_cmd_bits_isWr,
  output [25:0]  io_dram_cmd_bits_tag_uid,
  output [5:0]   io_dram_cmd_bits_tag_streamId,
  input          io_dram_wdata_ready,
  output         io_dram_wdata_valid,
  output [31:0]  io_dram_wdata_bits_wdata_0,
  output [31:0]  io_dram_wdata_bits_wdata_1,
  output [31:0]  io_dram_wdata_bits_wdata_2,
  output [31:0]  io_dram_wdata_bits_wdata_3,
  output [31:0]  io_dram_wdata_bits_wdata_4,
  output [31:0]  io_dram_wdata_bits_wdata_5,
  output [31:0]  io_dram_wdata_bits_wdata_6,
  output [31:0]  io_dram_wdata_bits_wdata_7,
  output [31:0]  io_dram_wdata_bits_wdata_8,
  output [31:0]  io_dram_wdata_bits_wdata_9,
  output [31:0]  io_dram_wdata_bits_wdata_10,
  output [31:0]  io_dram_wdata_bits_wdata_11,
  output [31:0]  io_dram_wdata_bits_wdata_12,
  output [31:0]  io_dram_wdata_bits_wdata_13,
  output [31:0]  io_dram_wdata_bits_wdata_14,
  output [31:0]  io_dram_wdata_bits_wdata_15,
  output         io_dram_wdata_bits_wstrb_0,
  output         io_dram_wdata_bits_wstrb_1,
  output         io_dram_wdata_bits_wstrb_2,
  output         io_dram_wdata_bits_wstrb_3,
  output         io_dram_wdata_bits_wstrb_4,
  output         io_dram_wdata_bits_wstrb_5,
  output         io_dram_wdata_bits_wstrb_6,
  output         io_dram_wdata_bits_wstrb_7,
  output         io_dram_wdata_bits_wstrb_8,
  output         io_dram_wdata_bits_wstrb_9,
  output         io_dram_wdata_bits_wstrb_10,
  output         io_dram_wdata_bits_wstrb_11,
  output         io_dram_wdata_bits_wstrb_12,
  output         io_dram_wdata_bits_wstrb_13,
  output         io_dram_wdata_bits_wstrb_14,
  output         io_dram_wdata_bits_wstrb_15,
  output         io_dram_wdata_bits_wstrb_16,
  output         io_dram_wdata_bits_wstrb_17,
  output         io_dram_wdata_bits_wstrb_18,
  output         io_dram_wdata_bits_wstrb_19,
  output         io_dram_wdata_bits_wstrb_20,
  output         io_dram_wdata_bits_wstrb_21,
  output         io_dram_wdata_bits_wstrb_22,
  output         io_dram_wdata_bits_wstrb_23,
  output         io_dram_wdata_bits_wstrb_24,
  output         io_dram_wdata_bits_wstrb_25,
  output         io_dram_wdata_bits_wstrb_26,
  output         io_dram_wdata_bits_wstrb_27,
  output         io_dram_wdata_bits_wstrb_28,
  output         io_dram_wdata_bits_wstrb_29,
  output         io_dram_wdata_bits_wstrb_30,
  output         io_dram_wdata_bits_wstrb_31,
  output         io_dram_wdata_bits_wstrb_32,
  output         io_dram_wdata_bits_wstrb_33,
  output         io_dram_wdata_bits_wstrb_34,
  output         io_dram_wdata_bits_wstrb_35,
  output         io_dram_wdata_bits_wstrb_36,
  output         io_dram_wdata_bits_wstrb_37,
  output         io_dram_wdata_bits_wstrb_38,
  output         io_dram_wdata_bits_wstrb_39,
  output         io_dram_wdata_bits_wstrb_40,
  output         io_dram_wdata_bits_wstrb_41,
  output         io_dram_wdata_bits_wstrb_42,
  output         io_dram_wdata_bits_wstrb_43,
  output         io_dram_wdata_bits_wstrb_44,
  output         io_dram_wdata_bits_wstrb_45,
  output         io_dram_wdata_bits_wstrb_46,
  output         io_dram_wdata_bits_wstrb_47,
  output         io_dram_wdata_bits_wstrb_48,
  output         io_dram_wdata_bits_wstrb_49,
  output         io_dram_wdata_bits_wstrb_50,
  output         io_dram_wdata_bits_wstrb_51,
  output         io_dram_wdata_bits_wstrb_52,
  output         io_dram_wdata_bits_wstrb_53,
  output         io_dram_wdata_bits_wstrb_54,
  output         io_dram_wdata_bits_wstrb_55,
  output         io_dram_wdata_bits_wstrb_56,
  output         io_dram_wdata_bits_wstrb_57,
  output         io_dram_wdata_bits_wstrb_58,
  output         io_dram_wdata_bits_wstrb_59,
  output         io_dram_wdata_bits_wstrb_60,
  output         io_dram_wdata_bits_wstrb_61,
  output         io_dram_wdata_bits_wstrb_62,
  output         io_dram_wdata_bits_wstrb_63,
  output         io_dram_rresp_ready,
  input          io_dram_rresp_valid,
  input  [31:0]  io_dram_rresp_bits_rdata_0,
  input  [31:0]  io_dram_rresp_bits_rdata_1,
  input  [31:0]  io_dram_rresp_bits_rdata_2,
  input  [31:0]  io_dram_rresp_bits_rdata_3,
  input  [31:0]  io_dram_rresp_bits_rdata_4,
  input  [31:0]  io_dram_rresp_bits_rdata_5,
  input  [31:0]  io_dram_rresp_bits_rdata_6,
  input  [31:0]  io_dram_rresp_bits_rdata_7,
  input  [31:0]  io_dram_rresp_bits_rdata_8,
  input  [31:0]  io_dram_rresp_bits_rdata_9,
  input  [31:0]  io_dram_rresp_bits_rdata_10,
  input  [31:0]  io_dram_rresp_bits_rdata_11,
  input  [31:0]  io_dram_rresp_bits_rdata_12,
  input  [31:0]  io_dram_rresp_bits_rdata_13,
  input  [31:0]  io_dram_rresp_bits_rdata_14,
  input  [31:0]  io_dram_rresp_bits_rdata_15,
  input  [5:0]   io_dram_rresp_bits_tag_streamId,
  output         io_dram_wresp_ready,
  input          io_dram_wresp_valid,
  input  [5:0]   io_dram_wresp_bits_tag_streamId,
  output [31:0]  io_debugSignals_0,
  output [31:0]  io_debugSignals_1,
  output [31:0]  io_debugSignals_2,
  output [31:0]  io_debugSignals_3,
  output [31:0]  io_debugSignals_4,
  output [31:0]  io_debugSignals_5,
  output [31:0]  io_debugSignals_6,
  output [31:0]  io_debugSignals_7,
  output [31:0]  io_debugSignals_8,
  output [31:0]  io_debugSignals_9,
  output [31:0]  io_debugSignals_10,
  output [31:0]  io_debugSignals_11,
  output [31:0]  io_debugSignals_12,
  output [31:0]  io_debugSignals_13,
  output [31:0]  io_debugSignals_14,
  output [31:0]  io_debugSignals_15,
  output [31:0]  io_debugSignals_16,
  output [31:0]  io_debugSignals_17,
  output [31:0]  io_debugSignals_18,
  output [31:0]  io_debugSignals_19,
  output [31:0]  io_debugSignals_20,
  output [31:0]  io_debugSignals_21,
  output [31:0]  io_debugSignals_22,
  output [31:0]  io_debugSignals_23,
  output [31:0]  io_debugSignals_24,
  output [31:0]  io_debugSignals_25,
  output [31:0]  io_debugSignals_26,
  output [31:0]  io_debugSignals_27,
  output [31:0]  io_debugSignals_28,
  output [31:0]  io_debugSignals_29,
  output [31:0]  io_debugSignals_30,
  output [31:0]  io_debugSignals_31,
  output [31:0]  io_debugSignals_32,
  output [31:0]  io_debugSignals_33,
  output [31:0]  io_debugSignals_34,
  output [31:0]  io_debugSignals_35,
  output [31:0]  io_debugSignals_36,
  output [31:0]  io_debugSignals_37,
  output [31:0]  io_debugSignals_38,
  output [31:0]  io_debugSignals_39,
  output [31:0]  io_debugSignals_40,
  output [31:0]  io_debugSignals_41,
  output [31:0]  io_debugSignals_42,
  output [31:0]  io_debugSignals_43,
  output [31:0]  io_debugSignals_44,
  output [31:0]  io_debugSignals_45,
  output [31:0]  io_debugSignals_46,
  output [31:0]  io_debugSignals_47,
  output [31:0]  io_debugSignals_48,
  output [31:0]  io_debugSignals_49,
  output [31:0]  io_debugSignals_50,
  output [31:0]  io_debugSignals_51,
  output [31:0]  io_debugSignals_52,
  output [31:0]  io_debugSignals_53,
  output [31:0]  io_debugSignals_54,
  output [31:0]  io_debugSignals_55,
  output [31:0]  io_debugSignals_56,
  output [31:0]  io_debugSignals_57,
  output [31:0]  io_debugSignals_58,
  output [31:0]  io_debugSignals_59,
  output [31:0]  io_debugSignals_60,
  output [31:0]  io_debugSignals_61,
  output [31:0]  io_debugSignals_62,
  output [31:0]  io_debugSignals_63,
  output [31:0]  io_debugSignals_64,
  output [31:0]  io_debugSignals_65,
  output [31:0]  io_debugSignals_66,
  output [31:0]  io_debugSignals_67,
  output [31:0]  io_debugSignals_68,
  output [31:0]  io_debugSignals_69,
  output [31:0]  io_debugSignals_70,
  output [31:0]  io_debugSignals_71,
  output [31:0]  io_debugSignals_72,
  output [31:0]  io_debugSignals_73,
  output [31:0]  io_debugSignals_74,
  output [31:0]  io_debugSignals_75,
  output [31:0]  io_debugSignals_76,
  output [31:0]  io_debugSignals_77,
  output [31:0]  io_debugSignals_78,
  output [31:0]  io_debugSignals_79,
  output [31:0]  io_debugSignals_80,
  output [31:0]  io_debugSignals_81,
  output [31:0]  io_debugSignals_82,
  output [31:0]  io_debugSignals_83,
  output [31:0]  io_debugSignals_84,
  output [31:0]  io_debugSignals_85,
  output [31:0]  io_debugSignals_86,
  output [31:0]  io_debugSignals_87,
  output [31:0]  io_debugSignals_88,
  output [31:0]  io_debugSignals_89,
  output [31:0]  io_debugSignals_90,
  output [31:0]  io_debugSignals_91,
  output [31:0]  io_debugSignals_92,
  output [31:0]  io_debugSignals_93,
  output [31:0]  io_debugSignals_94,
  output [31:0]  io_debugSignals_95,
  output [31:0]  io_debugSignals_96,
  output [31:0]  io_debugSignals_97,
  output [31:0]  io_debugSignals_98,
  output [31:0]  io_debugSignals_99,
  output [31:0]  io_debugSignals_100,
  output [31:0]  io_debugSignals_101,
  output [31:0]  io_debugSignals_102,
  output [31:0]  io_debugSignals_103,
  output [31:0]  io_debugSignals_104,
  output [31:0]  io_debugSignals_105,
  output [31:0]  io_debugSignals_106,
  output [31:0]  io_debugSignals_107,
  input  [63:0]  io_TOP_AXI_AWADDR,
  input  [7:0]   io_TOP_AXI_AWLEN,
  input          io_TOP_AXI_AWVALID,
  input          io_TOP_AXI_AWREADY,
  input          io_TOP_AXI_ARID,
  input  [63:0]  io_TOP_AXI_ARADDR,
  input  [7:0]   io_TOP_AXI_ARLEN,
  input  [2:0]   io_TOP_AXI_ARSIZE,
  input  [1:0]   io_TOP_AXI_ARBURST,
  input          io_TOP_AXI_ARVALID,
  input          io_TOP_AXI_ARREADY,
  input  [511:0] io_TOP_AXI_WDATA,
  input  [63:0]  io_TOP_AXI_WSTRB,
  input          io_TOP_AXI_WVALID,
  input          io_TOP_AXI_WREADY,
  input          io_TOP_AXI_RVALID,
  input          io_TOP_AXI_RREADY,
  input          io_TOP_AXI_BVALID,
  input          io_TOP_AXI_BREADY,
  input  [63:0]  io_DWIDTH_AXI_AWADDR,
  input  [7:0]   io_DWIDTH_AXI_AWLEN,
  input          io_DWIDTH_AXI_AWVALID,
  input          io_DWIDTH_AXI_AWREADY,
  input  [63:0]  io_DWIDTH_AXI_ARADDR,
  input  [7:0]   io_DWIDTH_AXI_ARLEN,
  input  [2:0]   io_DWIDTH_AXI_ARSIZE,
  input  [1:0]   io_DWIDTH_AXI_ARBURST,
  input          io_DWIDTH_AXI_ARVALID,
  input          io_DWIDTH_AXI_ARREADY,
  input  [511:0] io_DWIDTH_AXI_WDATA,
  input  [63:0]  io_DWIDTH_AXI_WSTRB,
  input          io_DWIDTH_AXI_WVALID,
  input          io_DWIDTH_AXI_WREADY,
  input          io_DWIDTH_AXI_RVALID,
  input          io_DWIDTH_AXI_RREADY,
  input          io_DWIDTH_AXI_BVALID,
  input          io_DWIDTH_AXI_BREADY
);
  wire  cmdArbiter_clock;
  wire  cmdArbiter_reset;
  wire [63:0] cmdArbiter_io_fifo_0_enq_0_addr;
  wire  cmdArbiter_io_fifo_0_enq_0_isWr;
  wire [15:0] cmdArbiter_io_fifo_0_enq_0_size;
  wire  cmdArbiter_io_fifo_0_enqVld;
  wire [63:0] cmdArbiter_io_fifo_0_deq_0_addr;
  wire  cmdArbiter_io_fifo_0_deq_0_isWr;
  wire [15:0] cmdArbiter_io_fifo_0_deq_0_size;
  wire  cmdArbiter_io_fifo_0_deqVld;
  wire  cmdArbiter_io_fifo_0_full;
  wire  cmdArbiter_io_fifo_0_empty;
  wire  cmdArbiter_io_fifo_0_almostEmpty;
  wire [63:0] cmdArbiter_io_fifo_1_deq_0_addr;
  wire  cmdArbiter_io_fifo_1_deq_0_isWr;
  wire [15:0] cmdArbiter_io_fifo_1_deq_0_size;
  wire  cmdArbiter_io_fifo_1_deqVld;
  wire  cmdArbiter_io_fifo_1_empty;
  wire [63:0] cmdArbiter_io_enq_0_0_addr;
  wire  cmdArbiter_io_enq_0_0_isWr;
  wire [15:0] cmdArbiter_io_enq_0_0_size;
  wire  cmdArbiter_io_enqVld_0;
  wire  cmdArbiter_io_full_0;
  wire [63:0] cmdArbiter_io_deq_0_addr;
  wire  cmdArbiter_io_deq_0_isWr;
  wire [15:0] cmdArbiter_io_deq_0_size;
  wire  cmdArbiter_io_deqVld;
  wire  cmdArbiter_io_deqReady;
  wire  cmdArbiter_io_empty;
  wire  cmdArbiter_io_tag;
  wire  cmdFifos_0_clock;
  wire  cmdFifos_0_reset;
  wire [63:0] cmdFifos_0_io_enq_0_addr;
  wire  cmdFifos_0_io_enq_0_isWr;
  wire [15:0] cmdFifos_0_io_enq_0_size;
  wire  cmdFifos_0_io_enqVld;
  wire [63:0] cmdFifos_0_io_deq_0_addr;
  wire  cmdFifos_0_io_deq_0_isWr;
  wire [15:0] cmdFifos_0_io_deq_0_size;
  wire  cmdFifos_0_io_deqVld;
  wire  cmdFifos_0_io_full;
  wire  cmdFifos_0_io_empty;
  wire  cmdFifos_0_io_almostEmpty;
  wire  cmdFifos_1_clock;
  wire  cmdFifos_1_reset;
  wire [63:0] cmdFifos_1_io_enq_0_addr;
  wire  cmdFifos_1_io_enq_0_isWr;
  wire [15:0] cmdFifos_1_io_enq_0_size;
  wire  cmdFifos_1_io_enqVld;
  wire [63:0] cmdFifos_1_io_deq_0_addr;
  wire  cmdFifos_1_io_deq_0_isWr;
  wire [15:0] cmdFifos_1_io_deq_0_size;
  wire  cmdFifos_1_io_deqVld;
  wire  cmdFifos_1_io_full;
  wire  cmdFifos_1_io_empty;
  wire  cmdFifos_1_io_almostEmpty;
  wire [31:0] _T_886;
  wire [63:0] _T_887;
  wire  FF_clock;
  wire  FF_reset;
  wire [63:0] FF_io_in;
  wire [63:0] FF_io_init;
  wire  FF_io_reset;
  wire [63:0] FF_io_out;
  wire  FF_io_enable;
  wire  sizeCounter_clock;
  wire  sizeCounter_reset;
  wire [15:0] sizeCounter_io_max;
  wire [15:0] sizeCounter_io_stride;
  wire [15:0] sizeCounter_io_out;
  wire  sizeCounter_io_last;
  wire  sizeCounter_io_reset;
  wire  sizeCounter_io_enable;
  wire  sizeCounter_io_done;
  wire  _T_891;
  wire [63:0] cmdAddr_bits;
  wire [63:0] _GEN_0;
  wire [64:0] _T_894;
  wire [63:0] _T_895;
  wire  _T_896;
  wire  _T_897;
  wire  cmdRead;
  wire  cmdWrite;
  wire  isSparseMux_io_ins_0;
  wire  isSparseMux_io_ins_1;
  wire  isSparseMux_io_sel;
  wire  isSparseMux_io_out;
  wire  burstCounter_clock;
  wire  burstCounter_reset;
  wire [15:0] burstCounter_io_max;
  wire [15:0] burstCounter_io_stride;
  wire [15:0] burstCounter_io_out;
  wire  burstCounter_io_last;
  wire  burstCounter_io_reset;
  wire  burstCounter_io_enable;
  wire  burstCounter_io_done;
  wire  burstTagCounter_clock;
  wire  burstTagCounter_reset;
  wire [9:0] burstTagCounter_io_out;
  wire  burstTagCounter_io_reset;
  wire  burstTagCounter_io_enable;
  wire  dramReadySeen;
  wire [15:0] _T_903;
  wire  cmdCooldown_clock;
  wire  cmdCooldown_reset;
  wire  cmdCooldown_io_in;
  wire  cmdCooldown_io_init;
  wire  cmdCooldown_io_reset;
  wire  cmdCooldown_io_out;
  wire  cmdCooldown_io_enable;
  wire  burstCounterDoneLatch_clock;
  wire  burstCounterDoneLatch_reset;
  wire  burstCounterDoneLatch_io_in;
  wire  burstCounterDoneLatch_io_init;
  wire  burstCounterDoneLatch_io_reset;
  wire  burstCounterDoneLatch_io_out;
  wire  burstCounterDoneLatch_io_enable;
  wire  sizeCounterDoneLatch_clock;
  wire  sizeCounterDoneLatch_reset;
  wire  sizeCounterDoneLatch_io_in;
  wire  sizeCounterDoneLatch_io_init;
  wire  sizeCounterDoneLatch_io_reset;
  wire  sizeCounterDoneLatch_io_out;
  wire  sizeCounterDoneLatch_io_enable;
  wire  _T_908;
  wire  rrespReadyMux_io_ins_0;
  wire  rrespReadyMux_io_out;
  wire  wdataMux_io_ins_0_valid;
  wire [31:0] wdataMux_io_ins_0_bits_wdata_0;
  wire [31:0] wdataMux_io_ins_0_bits_wdata_1;
  wire [31:0] wdataMux_io_ins_0_bits_wdata_2;
  wire [31:0] wdataMux_io_ins_0_bits_wdata_3;
  wire [31:0] wdataMux_io_ins_0_bits_wdata_4;
  wire [31:0] wdataMux_io_ins_0_bits_wdata_5;
  wire [31:0] wdataMux_io_ins_0_bits_wdata_6;
  wire [31:0] wdataMux_io_ins_0_bits_wdata_7;
  wire [31:0] wdataMux_io_ins_0_bits_wdata_8;
  wire [31:0] wdataMux_io_ins_0_bits_wdata_9;
  wire [31:0] wdataMux_io_ins_0_bits_wdata_10;
  wire [31:0] wdataMux_io_ins_0_bits_wdata_11;
  wire [31:0] wdataMux_io_ins_0_bits_wdata_12;
  wire [31:0] wdataMux_io_ins_0_bits_wdata_13;
  wire [31:0] wdataMux_io_ins_0_bits_wdata_14;
  wire [31:0] wdataMux_io_ins_0_bits_wdata_15;
  wire  wdataMux_io_ins_0_bits_wstrb_0;
  wire  wdataMux_io_ins_0_bits_wstrb_1;
  wire  wdataMux_io_ins_0_bits_wstrb_2;
  wire  wdataMux_io_ins_0_bits_wstrb_3;
  wire  wdataMux_io_ins_0_bits_wstrb_4;
  wire  wdataMux_io_ins_0_bits_wstrb_5;
  wire  wdataMux_io_ins_0_bits_wstrb_6;
  wire  wdataMux_io_ins_0_bits_wstrb_7;
  wire  wdataMux_io_ins_0_bits_wstrb_8;
  wire  wdataMux_io_ins_0_bits_wstrb_9;
  wire  wdataMux_io_ins_0_bits_wstrb_10;
  wire  wdataMux_io_ins_0_bits_wstrb_11;
  wire  wdataMux_io_ins_0_bits_wstrb_12;
  wire  wdataMux_io_ins_0_bits_wstrb_13;
  wire  wdataMux_io_ins_0_bits_wstrb_14;
  wire  wdataMux_io_ins_0_bits_wstrb_15;
  wire  wdataMux_io_ins_0_bits_wstrb_16;
  wire  wdataMux_io_ins_0_bits_wstrb_17;
  wire  wdataMux_io_ins_0_bits_wstrb_18;
  wire  wdataMux_io_ins_0_bits_wstrb_19;
  wire  wdataMux_io_ins_0_bits_wstrb_20;
  wire  wdataMux_io_ins_0_bits_wstrb_21;
  wire  wdataMux_io_ins_0_bits_wstrb_22;
  wire  wdataMux_io_ins_0_bits_wstrb_23;
  wire  wdataMux_io_ins_0_bits_wstrb_24;
  wire  wdataMux_io_ins_0_bits_wstrb_25;
  wire  wdataMux_io_ins_0_bits_wstrb_26;
  wire  wdataMux_io_ins_0_bits_wstrb_27;
  wire  wdataMux_io_ins_0_bits_wstrb_28;
  wire  wdataMux_io_ins_0_bits_wstrb_29;
  wire  wdataMux_io_ins_0_bits_wstrb_30;
  wire  wdataMux_io_ins_0_bits_wstrb_31;
  wire  wdataMux_io_ins_0_bits_wstrb_32;
  wire  wdataMux_io_ins_0_bits_wstrb_33;
  wire  wdataMux_io_ins_0_bits_wstrb_34;
  wire  wdataMux_io_ins_0_bits_wstrb_35;
  wire  wdataMux_io_ins_0_bits_wstrb_36;
  wire  wdataMux_io_ins_0_bits_wstrb_37;
  wire  wdataMux_io_ins_0_bits_wstrb_38;
  wire  wdataMux_io_ins_0_bits_wstrb_39;
  wire  wdataMux_io_ins_0_bits_wstrb_40;
  wire  wdataMux_io_ins_0_bits_wstrb_41;
  wire  wdataMux_io_ins_0_bits_wstrb_42;
  wire  wdataMux_io_ins_0_bits_wstrb_43;
  wire  wdataMux_io_ins_0_bits_wstrb_44;
  wire  wdataMux_io_ins_0_bits_wstrb_45;
  wire  wdataMux_io_ins_0_bits_wstrb_46;
  wire  wdataMux_io_ins_0_bits_wstrb_47;
  wire  wdataMux_io_ins_0_bits_wstrb_48;
  wire  wdataMux_io_ins_0_bits_wstrb_49;
  wire  wdataMux_io_ins_0_bits_wstrb_50;
  wire  wdataMux_io_ins_0_bits_wstrb_51;
  wire  wdataMux_io_ins_0_bits_wstrb_52;
  wire  wdataMux_io_ins_0_bits_wstrb_53;
  wire  wdataMux_io_ins_0_bits_wstrb_54;
  wire  wdataMux_io_ins_0_bits_wstrb_55;
  wire  wdataMux_io_ins_0_bits_wstrb_56;
  wire  wdataMux_io_ins_0_bits_wstrb_57;
  wire  wdataMux_io_ins_0_bits_wstrb_58;
  wire  wdataMux_io_ins_0_bits_wstrb_59;
  wire  wdataMux_io_ins_0_bits_wstrb_60;
  wire  wdataMux_io_ins_0_bits_wstrb_61;
  wire  wdataMux_io_ins_0_bits_wstrb_62;
  wire  wdataMux_io_ins_0_bits_wstrb_63;
  wire  wdataMux_io_out_valid;
  wire [31:0] wdataMux_io_out_bits_wdata_0;
  wire [31:0] wdataMux_io_out_bits_wdata_1;
  wire [31:0] wdataMux_io_out_bits_wdata_2;
  wire [31:0] wdataMux_io_out_bits_wdata_3;
  wire [31:0] wdataMux_io_out_bits_wdata_4;
  wire [31:0] wdataMux_io_out_bits_wdata_5;
  wire [31:0] wdataMux_io_out_bits_wdata_6;
  wire [31:0] wdataMux_io_out_bits_wdata_7;
  wire [31:0] wdataMux_io_out_bits_wdata_8;
  wire [31:0] wdataMux_io_out_bits_wdata_9;
  wire [31:0] wdataMux_io_out_bits_wdata_10;
  wire [31:0] wdataMux_io_out_bits_wdata_11;
  wire [31:0] wdataMux_io_out_bits_wdata_12;
  wire [31:0] wdataMux_io_out_bits_wdata_13;
  wire [31:0] wdataMux_io_out_bits_wdata_14;
  wire [31:0] wdataMux_io_out_bits_wdata_15;
  wire  wdataMux_io_out_bits_wstrb_0;
  wire  wdataMux_io_out_bits_wstrb_1;
  wire  wdataMux_io_out_bits_wstrb_2;
  wire  wdataMux_io_out_bits_wstrb_3;
  wire  wdataMux_io_out_bits_wstrb_4;
  wire  wdataMux_io_out_bits_wstrb_5;
  wire  wdataMux_io_out_bits_wstrb_6;
  wire  wdataMux_io_out_bits_wstrb_7;
  wire  wdataMux_io_out_bits_wstrb_8;
  wire  wdataMux_io_out_bits_wstrb_9;
  wire  wdataMux_io_out_bits_wstrb_10;
  wire  wdataMux_io_out_bits_wstrb_11;
  wire  wdataMux_io_out_bits_wstrb_12;
  wire  wdataMux_io_out_bits_wstrb_13;
  wire  wdataMux_io_out_bits_wstrb_14;
  wire  wdataMux_io_out_bits_wstrb_15;
  wire  wdataMux_io_out_bits_wstrb_16;
  wire  wdataMux_io_out_bits_wstrb_17;
  wire  wdataMux_io_out_bits_wstrb_18;
  wire  wdataMux_io_out_bits_wstrb_19;
  wire  wdataMux_io_out_bits_wstrb_20;
  wire  wdataMux_io_out_bits_wstrb_21;
  wire  wdataMux_io_out_bits_wstrb_22;
  wire  wdataMux_io_out_bits_wstrb_23;
  wire  wdataMux_io_out_bits_wstrb_24;
  wire  wdataMux_io_out_bits_wstrb_25;
  wire  wdataMux_io_out_bits_wstrb_26;
  wire  wdataMux_io_out_bits_wstrb_27;
  wire  wdataMux_io_out_bits_wstrb_28;
  wire  wdataMux_io_out_bits_wstrb_29;
  wire  wdataMux_io_out_bits_wstrb_30;
  wire  wdataMux_io_out_bits_wstrb_31;
  wire  wdataMux_io_out_bits_wstrb_32;
  wire  wdataMux_io_out_bits_wstrb_33;
  wire  wdataMux_io_out_bits_wstrb_34;
  wire  wdataMux_io_out_bits_wstrb_35;
  wire  wdataMux_io_out_bits_wstrb_36;
  wire  wdataMux_io_out_bits_wstrb_37;
  wire  wdataMux_io_out_bits_wstrb_38;
  wire  wdataMux_io_out_bits_wstrb_39;
  wire  wdataMux_io_out_bits_wstrb_40;
  wire  wdataMux_io_out_bits_wstrb_41;
  wire  wdataMux_io_out_bits_wstrb_42;
  wire  wdataMux_io_out_bits_wstrb_43;
  wire  wdataMux_io_out_bits_wstrb_44;
  wire  wdataMux_io_out_bits_wstrb_45;
  wire  wdataMux_io_out_bits_wstrb_46;
  wire  wdataMux_io_out_bits_wstrb_47;
  wire  wdataMux_io_out_bits_wstrb_48;
  wire  wdataMux_io_out_bits_wstrb_49;
  wire  wdataMux_io_out_bits_wstrb_50;
  wire  wdataMux_io_out_bits_wstrb_51;
  wire  wdataMux_io_out_bits_wstrb_52;
  wire  wdataMux_io_out_bits_wstrb_53;
  wire  wdataMux_io_out_bits_wstrb_54;
  wire  wdataMux_io_out_bits_wstrb_55;
  wire  wdataMux_io_out_bits_wstrb_56;
  wire  wdataMux_io_out_bits_wstrb_57;
  wire  wdataMux_io_out_bits_wstrb_58;
  wire  wdataMux_io_out_bits_wstrb_59;
  wire  wdataMux_io_out_bits_wstrb_60;
  wire  wdataMux_io_out_bits_wstrb_61;
  wire  wdataMux_io_out_bits_wstrb_62;
  wire  wdataMux_io_out_bits_wstrb_63;
  wire  cmdDeqValidMux_io_ins_0;
  wire  cmdDeqValidMux_io_ins_1;
  wire  cmdDeqValidMux_io_sel;
  wire  cmdDeqValidMux_io_out;
  wire  dramCmdMux_io_ins_0_valid;
  wire [63:0] dramCmdMux_io_ins_0_bits_addr;
  wire [31:0] dramCmdMux_io_ins_0_bits_size;
  wire  dramCmdMux_io_ins_0_bits_isWr;
  wire [25:0] dramCmdMux_io_ins_0_bits_tag_uid;
  wire [5:0] dramCmdMux_io_ins_0_bits_tag_streamId;
  wire  dramCmdMux_io_ins_1_valid;
  wire [63:0] dramCmdMux_io_ins_1_bits_addr;
  wire [31:0] dramCmdMux_io_ins_1_bits_size;
  wire  dramCmdMux_io_ins_1_bits_isWr;
  wire [25:0] dramCmdMux_io_ins_1_bits_tag_uid;
  wire [5:0] dramCmdMux_io_ins_1_bits_tag_streamId;
  wire  dramCmdMux_io_sel;
  wire  dramCmdMux_io_out_valid;
  wire [63:0] dramCmdMux_io_out_bits_addr;
  wire [31:0] dramCmdMux_io_out_bits_size;
  wire  dramCmdMux_io_out_bits_isWr;
  wire [25:0] dramCmdMux_io_out_bits_tag_uid;
  wire [5:0] dramCmdMux_io_out_bits_tag_streamId;
  wire [57:0] _T_931;
  wire [63:0] _T_933;
  wire [5:0] _T_935_streamId;
  wire [15:0] _T_937_bits;
  wire [16:0] _T_938;
  wire [16:0] _T_939;
  wire [15:0] _T_940;
  wire [15:0] _T_942;
  wire [15:0] _T_943;
  wire [9:0] _T_944;
  wire [5:0] _T_945;
  wire  _T_947;
  wire [9:0] _GEN_2;
  wire [10:0] _T_948;
  wire [9:0] _T_949;
  wire  _T_950;
  wire  _T_951;
  wire  FF_1_clock;
  wire  FF_1_reset;
  wire [5:0] FF_1_io_in;
  wire [5:0] FF_1_io_out;
  wire  FF_1_io_enable;
  wire  FF_2_clock;
  wire  FF_2_reset;
  wire [63:0] FF_2_io_in;
  wire [63:0] FF_2_io_init;
  wire  FF_2_io_reset;
  wire [63:0] FF_2_io_out;
  wire  FF_2_io_enable;
  wire  FF_3_clock;
  wire  FF_3_reset;
  wire [31:0] FF_3_io_in;
  wire [31:0] FF_3_io_out;
  wire  FF_3_io_enable;
  wire [5:0] _T_969_streamId;
  wire [15:0] _T_971_bits;
  wire [9:0] _T_978;
  wire [5:0] _T_979;
  wire  _T_981;
  wire [9:0] _GEN_3;
  wire [10:0] _T_982;
  wire [9:0] _T_983;
  wire  FF_4_clock;
  wire  FF_4_reset;
  wire  FF_4_io_in;
  wire  FF_4_io_init;
  wire  FF_4_io_reset;
  wire  FF_4_io_out;
  wire  FF_4_io_enable;
  wire  FF_5_clock;
  wire  FF_5_reset;
  wire [15:0] FF_5_io_in;
  wire [15:0] FF_5_io_out;
  wire  FF_5_io_enable;
  wire  wrespReadyMux_io_ins_0;
  wire  wrespReadyMux_io_out;
  wire  gatherLoadIssueMux_io_ins_0;
  wire  gatherLoadIssueMux_io_ins_1;
  wire  gatherLoadIssueMux_io_sel;
  wire  gatherLoadIssueMux_io_out;
  wire  gatherLoadIssue_clock;
  wire  gatherLoadIssue_reset;
  wire [63:0] gatherLoadIssue_io_out;
  wire  gatherLoadIssue_io_reset;
  wire  gatherLoadIssue_io_enable;
  wire  gatherLoadSkipMux_io_ins_0;
  wire  gatherLoadSkipMux_io_ins_1;
  wire  gatherLoadSkipMux_io_sel;
  wire  gatherLoadSkipMux_io_out;
  wire  gatherLoadSkip_clock;
  wire  gatherLoadSkip_reset;
  wire [63:0] gatherLoadSkip_io_out;
  wire  gatherLoadSkip_io_reset;
  wire  gatherLoadSkip_io_enable;
  wire  scatterLoadIssueMux_io_ins_0;
  wire  scatterLoadIssueMux_io_ins_1;
  wire  scatterLoadIssueMux_io_sel;
  wire  scatterLoadIssueMux_io_out;
  wire  scatterLoadIssue_clock;
  wire  scatterLoadIssue_reset;
  wire [63:0] scatterLoadIssue_io_out;
  wire  scatterLoadIssue_io_reset;
  wire  scatterLoadIssue_io_enable;
  wire  scatterLoadSkipMux_io_ins_0;
  wire  scatterLoadSkipMux_io_ins_1;
  wire  scatterLoadSkipMux_io_sel;
  wire  scatterLoadSkipMux_io_out;
  wire  scatterLoadSkip_clock;
  wire  scatterLoadSkip_reset;
  wire [63:0] scatterLoadSkip_io_out;
  wire  scatterLoadSkip_io_reset;
  wire  scatterLoadSkip_io_enable;
  wire  scatterStoreIssueMux_io_ins_0;
  wire  scatterStoreIssueMux_io_ins_1;
  wire  scatterStoreIssueMux_io_sel;
  wire  scatterStoreIssueMux_io_out;
  wire  scatterStoreIssue_clock;
  wire  scatterStoreIssue_reset;
  wire [63:0] scatterStoreIssue_io_out;
  wire  scatterStoreIssue_io_reset;
  wire  scatterStoreIssue_io_enable;
  wire  scatterStoreSkipMux_io_ins_0;
  wire  scatterStoreSkipMux_io_ins_1;
  wire  scatterStoreSkipMux_io_sel;
  wire  scatterStoreSkipMux_io_out;
  wire  scatterStoreSkip_clock;
  wire  scatterStoreSkip_reset;
  wire [63:0] scatterStoreSkip_io_out;
  wire  scatterStoreSkip_io_reset;
  wire  scatterStoreSkip_io_enable;
  wire  denseLoadBuffers_0_clock;
  wire  denseLoadBuffers_0_reset;
  wire [31:0] denseLoadBuffers_0_io_enq_0;
  wire [31:0] denseLoadBuffers_0_io_enq_1;
  wire [31:0] denseLoadBuffers_0_io_enq_2;
  wire [31:0] denseLoadBuffers_0_io_enq_3;
  wire [31:0] denseLoadBuffers_0_io_enq_4;
  wire [31:0] denseLoadBuffers_0_io_enq_5;
  wire [31:0] denseLoadBuffers_0_io_enq_6;
  wire [31:0] denseLoadBuffers_0_io_enq_7;
  wire [31:0] denseLoadBuffers_0_io_enq_8;
  wire [31:0] denseLoadBuffers_0_io_enq_9;
  wire [31:0] denseLoadBuffers_0_io_enq_10;
  wire [31:0] denseLoadBuffers_0_io_enq_11;
  wire [31:0] denseLoadBuffers_0_io_enq_12;
  wire [31:0] denseLoadBuffers_0_io_enq_13;
  wire [31:0] denseLoadBuffers_0_io_enq_14;
  wire [31:0] denseLoadBuffers_0_io_enq_15;
  wire  denseLoadBuffers_0_io_enqVld;
  wire [31:0] denseLoadBuffers_0_io_deq_0;
  wire  denseLoadBuffers_0_io_deqVld;
  wire  denseLoadBuffers_0_io_full;
  wire  denseLoadBuffers_0_io_empty;
  wire  denseLoadBuffers_0_io_almostEmpty;
  wire  denseLoadBuffers_0_io_almostFull;
  wire  _T_1027;
  wire  _T_1028;
  wire  _T_1029;
  wire  _T_1031;
  wire  Counter_clock;
  wire  Counter_reset;
  wire [63:0] Counter_io_out;
  wire  Counter_io_reset;
  wire  Counter_io_enable;
  wire  Counter_1_clock;
  wire  Counter_1_reset;
  wire [63:0] Counter_1_io_out;
  wire  Counter_1_io_reset;
  wire  Counter_1_io_enable;
  wire  Counter_2_clock;
  wire  Counter_2_reset;
  wire [63:0] Counter_2_io_out;
  wire  Counter_2_io_reset;
  wire  Counter_2_io_enable;
  wire  _T_1046;
  wire  Counter_3_clock;
  wire  Counter_3_reset;
  wire [63:0] Counter_3_io_out;
  wire  Counter_3_io_reset;
  wire  Counter_3_io_enable;
  wire  _T_1051;
  wire  Counter_4_clock;
  wire  Counter_4_reset;
  wire [63:0] Counter_4_io_out;
  wire  Counter_4_io_reset;
  wire  Counter_4_io_enable;
  wire  SRFF_clock;
  wire  SRFF_reset;
  wire  SRFF_io_input_set;
  wire  SRFF_io_input_reset;
  wire  SRFF_io_input_asyn_reset;
  wire  SRFF_io_output_data;
  wire  _T_1057;
  wire  SRFF_1_clock;
  wire  SRFF_1_reset;
  wire  SRFF_1_io_input_set;
  wire  SRFF_1_io_input_reset;
  wire  SRFF_1_io_input_asyn_reset;
  wire  SRFF_1_io_output_data;
  wire  _T_1064;
  wire  _T_1065;
  reg  _T_1068;
  reg [31:0] _RAND_0;
  wire  _T_1074;
  wire  _T_1075;
  wire  FF_6_clock;
  wire  FF_6_reset;
  wire [31:0] FF_6_io_in;
  wire [31:0] FF_6_io_out;
  wire  FF_6_io_enable;
  wire  _T_1079;
  wire  _T_1080;
  reg  _T_1083;
  reg [31:0] _RAND_1;
  wire  _T_1089;
  wire  _T_1090;
  wire [63:0] _T_1091;
  wire [95:0] _T_1092;
  wire [127:0] _T_1093;
  wire [159:0] _T_1094;
  wire [191:0] _T_1095;
  wire [223:0] _T_1096;
  wire [255:0] _T_1097;
  wire [287:0] _T_1098;
  wire [319:0] _T_1099;
  wire [351:0] _T_1100;
  wire [383:0] _T_1101;
  wire [415:0] _T_1102;
  wire [447:0] _T_1103;
  wire [479:0] _T_1104;
  wire [511:0] _T_1105;
  wire  FF_7_clock;
  wire  FF_7_reset;
  wire [511:0] FF_7_io_in;
  wire [511:0] FF_7_io_out;
  wire  FF_7_io_enable;
  wire  denseStoreBuffers_0_clock;
  wire  denseStoreBuffers_0_reset;
  wire  denseStoreBuffers_0_io_enqVld;
  wire [31:0] denseStoreBuffers_0_io_deq_0;
  wire [31:0] denseStoreBuffers_0_io_deq_1;
  wire [31:0] denseStoreBuffers_0_io_deq_2;
  wire [31:0] denseStoreBuffers_0_io_deq_3;
  wire [31:0] denseStoreBuffers_0_io_deq_4;
  wire [31:0] denseStoreBuffers_0_io_deq_5;
  wire [31:0] denseStoreBuffers_0_io_deq_6;
  wire [31:0] denseStoreBuffers_0_io_deq_7;
  wire [31:0] denseStoreBuffers_0_io_deq_8;
  wire [31:0] denseStoreBuffers_0_io_deq_9;
  wire [31:0] denseStoreBuffers_0_io_deq_10;
  wire [31:0] denseStoreBuffers_0_io_deq_11;
  wire [31:0] denseStoreBuffers_0_io_deq_12;
  wire [31:0] denseStoreBuffers_0_io_deq_13;
  wire [31:0] denseStoreBuffers_0_io_deq_14;
  wire [31:0] denseStoreBuffers_0_io_deq_15;
  wire [63:0] denseStoreBuffers_0_io_deqStrb;
  wire  denseStoreBuffers_0_io_deqVld;
  wire  denseStoreBuffers_0_io_full;
  wire  denseStoreBuffers_0_io_empty;
  wire  denseStoreBuffers_0_io_almostEmpty;
  wire  denseStoreBuffers_0_io_almostFull;
  wire  _T_1109;
  wire  _T_1110;
  wire  _T_1111;
  wire  _T_1112;
  wire  _T_1114;
  wire  _T_1115;
  wire  _T_1116;
  wire  _T_1118;
  wire  _T_1119;
  wire  _T_1120;
  wire  _T_1121;
  wire  _T_1122;
  wire  _T_1123;
  wire  _T_1127;
  wire  _T_1129;
  wire  _T_1130;
  wire  _T_1131;
  wire  _T_1132;
  wire  _T_1133;
  wire  _T_1134;
  wire  _T_1135;
  wire  _T_1136;
  wire  _T_1137;
  wire  _T_1138;
  wire  _T_1139;
  wire  _T_1140;
  wire  _T_1141;
  wire  _T_1142;
  wire  _T_1143;
  wire  _T_1144;
  wire  _T_1145;
  wire  _T_1146;
  wire  _T_1147;
  wire  _T_1148;
  wire  _T_1149;
  wire  _T_1150;
  wire  _T_1151;
  wire  _T_1152;
  wire  _T_1153;
  wire  _T_1154;
  wire  _T_1155;
  wire  _T_1156;
  wire  _T_1157;
  wire  _T_1158;
  wire  _T_1159;
  wire  _T_1160;
  wire  _T_1161;
  wire  _T_1162;
  wire  _T_1163;
  wire  _T_1164;
  wire  _T_1165;
  wire  _T_1166;
  wire  _T_1167;
  wire  _T_1168;
  wire  _T_1169;
  wire  _T_1170;
  wire  _T_1171;
  wire  _T_1172;
  wire  _T_1173;
  wire  _T_1174;
  wire  _T_1175;
  wire  _T_1176;
  wire  _T_1177;
  wire  _T_1178;
  wire  _T_1179;
  wire  _T_1180;
  wire  _T_1181;
  wire  _T_1182;
  wire  _T_1183;
  wire  _T_1184;
  wire  _T_1185;
  wire  _T_1186;
  wire  _T_1187;
  wire  _T_1188;
  wire  _T_1189;
  wire  _T_1190;
  wire  _T_1191;
  wire  _T_1192;
  wire  _T_1193;
  wire  _T_1194;
  wire  Counter_5_clock;
  wire  Counter_5_reset;
  wire [15:0] Counter_5_io_max;
  wire [15:0] Counter_5_io_stride;
  wire [15:0] Counter_5_io_out;
  wire  Counter_5_io_last;
  wire  Counter_5_io_reset;
  wire  Counter_5_io_enable;
  wire  Counter_5_io_done;
  wire  FF_8_clock;
  wire  FF_8_reset;
  wire [15:0] FF_8_io_in;
  wire [15:0] FF_8_io_out;
  wire  FF_8_io_enable;
  wire  _T_1197;
  wire  _T_1202;
  wire  _T_1203;
  wire  FIFOCounter_clock;
  wire  FIFOCounter_reset;
  wire  FIFOCounter_io_enqVld;
  wire  FIFOCounter_io_full;
  wire  FIFOCounter_io_empty;
  wire  _T_1204;
  wire  _T_1205;
  wire  Counter_6_clock;
  wire  Counter_6_reset;
  wire [63:0] Counter_6_io_out;
  wire  Counter_6_io_reset;
  wire  Counter_6_io_enable;
  wire  Counter_7_clock;
  wire  Counter_7_reset;
  wire [63:0] Counter_7_io_out;
  wire  Counter_7_io_reset;
  wire  Counter_7_io_enable;
  wire  Counter_8_clock;
  wire  Counter_8_reset;
  wire [63:0] Counter_8_io_out;
  wire  Counter_8_io_reset;
  wire  Counter_8_io_enable;
  wire  burstCounterMaxLatch_clock;
  wire  burstCounterMaxLatch_reset;
  wire [31:0] burstCounterMaxLatch_io_in;
  wire [31:0] burstCounterMaxLatch_io_out;
  wire  burstCounterMaxLatch_io_enable;
  wire [31:0] burstCounterMax;
  wire  _T_1227;
  wire  _T_1229;
  wire [31:0] _T_1231;
  wire  _T_1233;
  wire  _T_1235;
  wire  dramReadyFF_clock;
  wire  dramReadyFF_reset;
  wire  dramReadyFF_io_in;
  wire  dramReadyFF_io_init;
  wire  dramReadyFF_io_reset;
  wire  dramReadyFF_io_out;
  wire  dramReadyFF_io_enable;
  wire  dramReadyFFEnabler;
  wire  _T_1243;
  wire  _T_1244;
  wire  _T_1246;
  wire  _T_1247;
  wire  _T_1249;
  wire  _T_1255;
  wire  _T_1256;
  wire  cycleCount_clock;
  wire  cycleCount_reset;
  wire [63:0] cycleCount_io_out;
  wire  cycleCount_io_reset;
  wire  cycleCount_io_enable;
  wire  _T_1261;
  wire  rdataEnqCount_clock;
  wire  rdataEnqCount_reset;
  wire [63:0] rdataEnqCount_io_out;
  wire  rdataEnqCount_io_reset;
  wire  rdataEnqCount_io_enable;
  wire  _T_1266;
  wire  _T_1267;
  wire  wdataCount_clock;
  wire  wdataCount_reset;
  wire [63:0] wdataCount_io_out;
  wire  wdataCount_io_reset;
  wire  wdataCount_io_enable;
  wire  _T_1272;
  wire  _T_1273;
  wire  Counter_9_clock;
  wire  Counter_9_reset;
  wire [63:0] Counter_9_io_out;
  wire  Counter_9_io_reset;
  wire  Counter_9_io_enable;
  wire  _T_1278;
  wire  _T_1279;
  wire  _T_1280;
  wire  _T_1281;
  wire  _T_1282;
  wire  Counter_10_clock;
  wire  Counter_10_reset;
  wire [63:0] Counter_10_io_out;
  wire  Counter_10_io_reset;
  wire  Counter_10_io_enable;
  wire  _T_1290;
  wire  Counter_11_clock;
  wire  Counter_11_reset;
  wire [63:0] Counter_11_io_out;
  wire  Counter_11_io_reset;
  wire  Counter_11_io_enable;
  wire  _T_1295;
  wire  Counter_12_clock;
  wire  Counter_12_reset;
  wire [63:0] Counter_12_io_out;
  wire  Counter_12_io_reset;
  wire  Counter_12_io_enable;
  wire  _T_1301;
  wire  Counter_13_clock;
  wire  Counter_13_reset;
  wire [63:0] Counter_13_io_out;
  wire  Counter_13_io_reset;
  wire  Counter_13_io_enable;
  wire  _T_1308;
  wire  _T_1309;
  wire  Counter_14_clock;
  wire  Counter_14_reset;
  wire [63:0] Counter_14_io_out;
  wire  Counter_14_io_reset;
  wire  Counter_14_io_enable;
  wire  _T_1316;
  wire  Counter_15_clock;
  wire  Counter_15_reset;
  wire [63:0] Counter_15_io_out;
  wire  Counter_15_io_reset;
  wire  Counter_15_io_enable;
  wire  Counter_16_clock;
  wire  Counter_16_reset;
  wire [63:0] Counter_16_io_out;
  wire  Counter_16_io_reset;
  wire  Counter_16_io_enable;
  wire  Counter_17_clock;
  wire  Counter_17_reset;
  wire [63:0] Counter_17_io_out;
  wire  Counter_17_io_reset;
  wire  Counter_17_io_enable;
  wire  _T_1335;
  wire  Counter_18_clock;
  wire  Counter_18_reset;
  wire [63:0] Counter_18_io_out;
  wire  Counter_18_io_reset;
  wire  Counter_18_io_enable;
  wire  Counter_19_clock;
  wire  Counter_19_reset;
  wire [63:0] Counter_19_io_out;
  wire  Counter_19_io_reset;
  wire  Counter_19_io_enable;
  wire  _T_1345;
  wire  _T_1346;
  wire  _T_1347;
  wire  Counter_20_clock;
  wire  Counter_20_reset;
  wire [63:0] Counter_20_io_out;
  wire  Counter_20_io_reset;
  wire  Counter_20_io_enable;
  wire  _T_1352;
  wire  _T_1353;
  wire  _T_1354;
  wire  Counter_21_clock;
  wire  Counter_21_reset;
  wire [63:0] Counter_21_io_out;
  wire  Counter_21_io_reset;
  wire  Counter_21_io_enable;
  wire  _T_1362;
  wire  Counter_22_clock;
  wire  Counter_22_reset;
  wire [63:0] Counter_22_io_out;
  wire  Counter_22_io_reset;
  wire  Counter_22_io_enable;
  wire  _T_1367;
  wire  Counter_23_clock;
  wire  Counter_23_reset;
  wire [63:0] Counter_23_io_out;
  wire  Counter_23_io_reset;
  wire  Counter_23_io_enable;
  wire  _T_1372;
  wire  _T_1373;
  wire  _T_1374;
  wire  Counter_24_clock;
  wire  Counter_24_reset;
  wire [63:0] Counter_24_io_out;
  wire  Counter_24_io_reset;
  wire  Counter_24_io_enable;
  wire  _T_1379;
  wire  _T_1380;
  wire  _T_1381;
  wire  Counter_25_clock;
  wire  Counter_25_reset;
  wire [63:0] Counter_25_io_out;
  wire  Counter_25_io_reset;
  wire  Counter_25_io_enable;
  wire  _T_1389;
  wire  Counter_26_clock;
  wire  Counter_26_reset;
  wire [63:0] Counter_26_io_out;
  wire  Counter_26_io_reset;
  wire  Counter_26_io_enable;
  wire  Counter_27_clock;
  wire  Counter_27_reset;
  wire [63:0] Counter_27_io_out;
  wire  Counter_27_io_reset;
  wire  Counter_27_io_enable;
  wire  Counter_28_clock;
  wire  Counter_28_reset;
  wire [63:0] Counter_28_io_out;
  wire  Counter_28_io_reset;
  wire  Counter_28_io_enable;
  wire  Counter_29_clock;
  wire  Counter_29_reset;
  wire [63:0] Counter_29_io_out;
  wire  Counter_29_io_reset;
  wire  Counter_29_io_enable;
  wire  Counter_30_clock;
  wire  Counter_30_reset;
  wire [63:0] Counter_30_io_out;
  wire  Counter_30_io_reset;
  wire  Counter_30_io_enable;
  wire  Counter_31_clock;
  wire  Counter_31_reset;
  wire [63:0] Counter_31_io_out;
  wire  Counter_31_io_reset;
  wire  Counter_31_io_enable;
  wire  Counter_32_clock;
  wire  Counter_32_reset;
  wire [63:0] Counter_32_io_out;
  wire  Counter_32_io_reset;
  wire  Counter_32_io_enable;
  wire  Counter_33_clock;
  wire  Counter_33_reset;
  wire [63:0] Counter_33_io_out;
  wire  Counter_33_io_reset;
  wire  Counter_33_io_enable;
  wire  _T_1425;
  wire  Counter_34_clock;
  wire  Counter_34_reset;
  wire [63:0] Counter_34_io_out;
  wire  Counter_34_io_reset;
  wire  Counter_34_io_enable;
  wire  FF_9_clock;
  wire  FF_9_reset;
  wire [5:0] FF_9_io_in;
  wire [5:0] FF_9_io_out;
  wire  FF_9_io_enable;
  wire  Counter_35_clock;
  wire  Counter_35_reset;
  wire [63:0] Counter_35_io_out;
  wire  Counter_35_io_reset;
  wire  Counter_35_io_enable;
  wire  Counter_36_clock;
  wire  Counter_36_reset;
  wire [63:0] Counter_36_io_out;
  wire  Counter_36_io_reset;
  wire  Counter_36_io_enable;
  wire  _T_1443;
  wire  Counter_37_clock;
  wire  Counter_37_reset;
  wire [63:0] Counter_37_io_out;
  wire  Counter_37_io_reset;
  wire  Counter_37_io_enable;
  wire  _T_1448;
  wire  Counter_38_clock;
  wire  Counter_38_reset;
  wire [63:0] Counter_38_io_out;
  wire  Counter_38_io_reset;
  wire  Counter_38_io_enable;
  wire  Counter_39_clock;
  wire  Counter_39_reset;
  wire [63:0] Counter_39_io_out;
  wire  Counter_39_io_reset;
  wire  Counter_39_io_enable;
  wire  Counter_40_clock;
  wire  Counter_40_reset;
  wire [63:0] Counter_40_io_out;
  wire  Counter_40_io_reset;
  wire  Counter_40_io_enable;
  wire  Counter_41_clock;
  wire  Counter_41_reset;
  wire [63:0] Counter_41_io_out;
  wire  Counter_41_io_reset;
  wire  Counter_41_io_enable;
  wire  Counter_42_clock;
  wire  Counter_42_reset;
  wire [63:0] Counter_42_io_out;
  wire  Counter_42_io_reset;
  wire  Counter_42_io_enable;
  wire  _T_1469;
  wire  Counter_43_clock;
  wire  Counter_43_reset;
  wire [63:0] Counter_43_io_out;
  wire  Counter_43_io_reset;
  wire  Counter_43_io_enable;
  wire  Counter_44_clock;
  wire  Counter_44_reset;
  wire [63:0] Counter_44_io_out;
  wire  Counter_44_io_reset;
  wire  Counter_44_io_enable;
  wire  _T_1480;
  wire  Counter_45_clock;
  wire  Counter_45_reset;
  wire [63:0] Counter_45_io_out;
  wire  Counter_45_io_reset;
  wire  Counter_45_io_enable;
  wire  _T_1486;
  wire  Counter_46_clock;
  wire  Counter_46_reset;
  wire [63:0] Counter_46_io_out;
  wire  Counter_46_io_reset;
  wire  Counter_46_io_enable;
  wire  Counter_47_clock;
  wire  Counter_47_reset;
  wire [63:0] Counter_47_io_out;
  wire  Counter_47_io_reset;
  wire  Counter_47_io_enable;
  wire  Counter_48_clock;
  wire  Counter_48_reset;
  wire [63:0] Counter_48_io_out;
  wire  Counter_48_io_reset;
  wire  Counter_48_io_enable;
  wire  _T_1499;
  wire  Counter_49_clock;
  wire  Counter_49_reset;
  wire [63:0] Counter_49_io_out;
  wire  Counter_49_io_reset;
  wire  Counter_49_io_enable;
  wire  Counter_50_clock;
  wire  Counter_50_reset;
  wire [63:0] Counter_50_io_out;
  wire  Counter_50_io_reset;
  wire  Counter_50_io_enable;
  wire  _T_1508;
  wire  Counter_51_clock;
  wire  Counter_51_reset;
  wire [63:0] Counter_51_io_out;
  wire  Counter_51_io_reset;
  wire  Counter_51_io_enable;
  wire  Counter_52_clock;
  wire  Counter_52_reset;
  wire [63:0] Counter_52_io_out;
  wire  Counter_52_io_reset;
  wire  Counter_52_io_enable;
  wire  _T_1517;
  wire  Counter_53_clock;
  wire  Counter_53_reset;
  wire [63:0] Counter_53_io_out;
  wire  Counter_53_io_reset;
  wire  Counter_53_io_enable;
  wire  Counter_54_clock;
  wire  Counter_54_reset;
  wire [63:0] Counter_54_io_out;
  wire  Counter_54_io_reset;
  wire  Counter_54_io_enable;
  wire  _T_1526;
  wire  Counter_55_clock;
  wire  Counter_55_reset;
  wire [63:0] Counter_55_io_out;
  wire  Counter_55_io_reset;
  wire  Counter_55_io_enable;
  wire  _T_1531;
  wire  _T_1532;
  wire  Counter_56_clock;
  wire  Counter_56_reset;
  wire [63:0] Counter_56_io_out;
  wire  Counter_56_io_reset;
  wire  Counter_56_io_enable;
  wire  Counter_57_clock;
  wire  Counter_57_reset;
  wire [63:0] Counter_57_io_out;
  wire  Counter_57_io_reset;
  wire  Counter_57_io_enable;
  wire  Counter_58_clock;
  wire  Counter_58_reset;
  wire [63:0] Counter_58_io_out;
  wire  Counter_58_io_reset;
  wire  Counter_58_io_enable;
  wire  _T_1546;
  wire  Counter_59_clock;
  wire  Counter_59_reset;
  wire [63:0] Counter_59_io_out;
  wire  Counter_59_io_reset;
  wire  Counter_59_io_enable;
  wire  _T_1551;
  wire  FF_10_clock;
  wire  FF_10_reset;
  wire [63:0] FF_10_io_in;
  wire [63:0] FF_10_io_init;
  wire  FF_10_io_reset;
  wire [63:0] FF_10_io_out;
  wire  FF_10_io_enable;
  wire  FF_11_clock;
  wire  FF_11_reset;
  wire [7:0] FF_11_io_in;
  wire [7:0] FF_11_io_out;
  wire  FF_11_io_enable;
  wire  FF_12_clock;
  wire  FF_12_reset;
  wire [2:0] FF_12_io_in;
  wire [2:0] FF_12_io_out;
  wire  FF_12_io_enable;
  wire  FF_13_clock;
  wire  FF_13_reset;
  wire  FF_13_io_in;
  wire  FF_13_io_init;
  wire  FF_13_io_reset;
  wire  FF_13_io_out;
  wire  FF_13_io_enable;
  wire  FF_14_clock;
  wire  FF_14_reset;
  wire [1:0] FF_14_io_in;
  wire [1:0] FF_14_io_out;
  wire  FF_14_io_enable;
  wire  _T_1571;
  wire  FF_15_clock;
  wire  FF_15_reset;
  wire [63:0] FF_15_io_in;
  wire [63:0] FF_15_io_init;
  wire  FF_15_io_reset;
  wire [63:0] FF_15_io_out;
  wire  FF_15_io_enable;
  wire  FF_16_clock;
  wire  FF_16_reset;
  wire [7:0] FF_16_io_in;
  wire [7:0] FF_16_io_out;
  wire  FF_16_io_enable;
  wire  _T_1579;
  wire  FF_17_clock;
  wire  FF_17_reset;
  wire [511:0] FF_17_io_in;
  wire [511:0] FF_17_io_out;
  wire  FF_17_io_enable;
  wire  FF_18_clock;
  wire  FF_18_reset;
  wire [63:0] FF_18_io_in;
  wire [63:0] FF_18_io_init;
  wire  FF_18_io_reset;
  wire [63:0] FF_18_io_out;
  wire  FF_18_io_enable;
  wire  _T_1589;
  wire  _T_1590;
  wire  FF_19_clock;
  wire  FF_19_reset;
  wire [511:0] FF_19_io_in;
  wire [511:0] FF_19_io_out;
  wire  FF_19_io_enable;
  wire  FF_20_clock;
  wire  FF_20_reset;
  wire [63:0] FF_20_io_in;
  wire [63:0] FF_20_io_init;
  wire  FF_20_io_reset;
  wire [63:0] FF_20_io_out;
  wire  FF_20_io_enable;
  wire  _T_1603;
  wire  _T_1604;
  wire  FF_21_clock;
  wire  FF_21_reset;
  wire [511:0] FF_21_io_in;
  wire [511:0] FF_21_io_out;
  wire  FF_21_io_enable;
  wire  FF_22_clock;
  wire  FF_22_reset;
  wire [63:0] FF_22_io_in;
  wire [63:0] FF_22_io_init;
  wire  FF_22_io_reset;
  wire [63:0] FF_22_io_out;
  wire  FF_22_io_enable;
  wire  Counter_60_clock;
  wire  Counter_60_reset;
  wire [63:0] Counter_60_io_out;
  wire  Counter_60_io_reset;
  wire  Counter_60_io_enable;
  wire  Counter_61_clock;
  wire  Counter_61_reset;
  wire [63:0] Counter_61_io_out;
  wire  Counter_61_io_reset;
  wire  Counter_61_io_enable;
  wire  _T_1623;
  wire  Counter_62_clock;
  wire  Counter_62_reset;
  wire [63:0] Counter_62_io_out;
  wire  Counter_62_io_reset;
  wire  Counter_62_io_enable;
  wire  Counter_63_clock;
  wire  Counter_63_reset;
  wire [63:0] Counter_63_io_out;
  wire  Counter_63_io_reset;
  wire  Counter_63_io_enable;
  wire  _T_1632;
  wire  Counter_64_clock;
  wire  Counter_64_reset;
  wire [63:0] Counter_64_io_out;
  wire  Counter_64_io_reset;
  wire  Counter_64_io_enable;
  wire  Counter_65_clock;
  wire  Counter_65_reset;
  wire [63:0] Counter_65_io_out;
  wire  Counter_65_io_reset;
  wire  Counter_65_io_enable;
  wire  _T_1641;
  wire  Counter_66_clock;
  wire  Counter_66_reset;
  wire [63:0] Counter_66_io_out;
  wire  Counter_66_io_reset;
  wire  Counter_66_io_enable;
  wire  Counter_67_clock;
  wire  Counter_67_reset;
  wire [63:0] Counter_67_io_out;
  wire  Counter_67_io_reset;
  wire  Counter_67_io_enable;
  wire  _T_1650;
  wire  Counter_68_clock;
  wire  Counter_68_reset;
  wire [63:0] Counter_68_io_out;
  wire  Counter_68_io_reset;
  wire  Counter_68_io_enable;
  wire  _T_1655;
  wire  _T_1656;
  wire  Counter_69_clock;
  wire  Counter_69_reset;
  wire [63:0] Counter_69_io_out;
  wire  Counter_69_io_reset;
  wire  Counter_69_io_enable;
  wire  Counter_70_clock;
  wire  Counter_70_reset;
  wire [63:0] Counter_70_io_out;
  wire  Counter_70_io_reset;
  wire  Counter_70_io_enable;
  wire  Counter_71_clock;
  wire  Counter_71_reset;
  wire [63:0] Counter_71_io_out;
  wire  Counter_71_io_reset;
  wire  Counter_71_io_enable;
  wire  _T_1670;
  wire  Counter_72_clock;
  wire  Counter_72_reset;
  wire [63:0] Counter_72_io_out;
  wire  Counter_72_io_reset;
  wire  Counter_72_io_enable;
  wire  _T_1675;
  wire  FF_23_clock;
  wire  FF_23_reset;
  wire [63:0] FF_23_io_in;
  wire [63:0] FF_23_io_init;
  wire  FF_23_io_reset;
  wire [63:0] FF_23_io_out;
  wire  FF_23_io_enable;
  wire  FF_24_clock;
  wire  FF_24_reset;
  wire [7:0] FF_24_io_in;
  wire [7:0] FF_24_io_out;
  wire  FF_24_io_enable;
  wire  FF_25_clock;
  wire  FF_25_reset;
  wire [2:0] FF_25_io_in;
  wire [2:0] FF_25_io_out;
  wire  FF_25_io_enable;
  wire  FF_26_clock;
  wire  FF_26_reset;
  wire [1:0] FF_26_io_in;
  wire [1:0] FF_26_io_out;
  wire  FF_26_io_enable;
  wire  _T_1691;
  wire  FF_27_clock;
  wire  FF_27_reset;
  wire [63:0] FF_27_io_in;
  wire [63:0] FF_27_io_init;
  wire  FF_27_io_reset;
  wire [63:0] FF_27_io_out;
  wire  FF_27_io_enable;
  wire  FF_28_clock;
  wire  FF_28_reset;
  wire [7:0] FF_28_io_in;
  wire [7:0] FF_28_io_out;
  wire  FF_28_io_enable;
  wire  _T_1699;
  wire  FF_29_clock;
  wire  FF_29_reset;
  wire [511:0] FF_29_io_in;
  wire [511:0] FF_29_io_out;
  wire  FF_29_io_enable;
  wire  FF_30_clock;
  wire  FF_30_reset;
  wire [63:0] FF_30_io_in;
  wire [63:0] FF_30_io_init;
  wire  FF_30_io_reset;
  wire [63:0] FF_30_io_out;
  wire  FF_30_io_enable;
  wire  _T_1710;
  wire  FF_31_clock;
  wire  FF_31_reset;
  wire [511:0] FF_31_io_in;
  wire [511:0] FF_31_io_out;
  wire  FF_31_io_enable;
  wire  FF_32_clock;
  wire  FF_32_reset;
  wire [63:0] FF_32_io_in;
  wire [63:0] FF_32_io_init;
  wire  FF_32_io_reset;
  wire [63:0] FF_32_io_out;
  wire  FF_32_io_enable;
  wire  _T_1724;
  wire  FF_33_clock;
  wire  FF_33_reset;
  wire [511:0] FF_33_io_in;
  wire [511:0] FF_33_io_out;
  wire  FF_33_io_enable;
  wire  FF_34_clock;
  wire  FF_34_reset;
  wire [63:0] FF_34_io_in;
  wire [63:0] FF_34_io_init;
  wire  FF_34_io_reset;
  wire [63:0] FF_34_io_out;
  wire  FF_34_io_enable;
  FIFOArbiter cmdArbiter (
    .clock(cmdArbiter_clock),
    .reset(cmdArbiter_reset),
    .io_fifo_0_enq_0_addr(cmdArbiter_io_fifo_0_enq_0_addr),
    .io_fifo_0_enq_0_isWr(cmdArbiter_io_fifo_0_enq_0_isWr),
    .io_fifo_0_enq_0_size(cmdArbiter_io_fifo_0_enq_0_size),
    .io_fifo_0_enqVld(cmdArbiter_io_fifo_0_enqVld),
    .io_fifo_0_deq_0_addr(cmdArbiter_io_fifo_0_deq_0_addr),
    .io_fifo_0_deq_0_isWr(cmdArbiter_io_fifo_0_deq_0_isWr),
    .io_fifo_0_deq_0_size(cmdArbiter_io_fifo_0_deq_0_size),
    .io_fifo_0_deqVld(cmdArbiter_io_fifo_0_deqVld),
    .io_fifo_0_full(cmdArbiter_io_fifo_0_full),
    .io_fifo_0_empty(cmdArbiter_io_fifo_0_empty),
    .io_fifo_0_almostEmpty(cmdArbiter_io_fifo_0_almostEmpty),
    .io_fifo_1_deq_0_addr(cmdArbiter_io_fifo_1_deq_0_addr),
    .io_fifo_1_deq_0_isWr(cmdArbiter_io_fifo_1_deq_0_isWr),
    .io_fifo_1_deq_0_size(cmdArbiter_io_fifo_1_deq_0_size),
    .io_fifo_1_deqVld(cmdArbiter_io_fifo_1_deqVld),
    .io_fifo_1_empty(cmdArbiter_io_fifo_1_empty),
    .io_enq_0_0_addr(cmdArbiter_io_enq_0_0_addr),
    .io_enq_0_0_isWr(cmdArbiter_io_enq_0_0_isWr),
    .io_enq_0_0_size(cmdArbiter_io_enq_0_0_size),
    .io_enqVld_0(cmdArbiter_io_enqVld_0),
    .io_full_0(cmdArbiter_io_full_0),
    .io_deq_0_addr(cmdArbiter_io_deq_0_addr),
    .io_deq_0_isWr(cmdArbiter_io_deq_0_isWr),
    .io_deq_0_size(cmdArbiter_io_deq_0_size),
    .io_deqVld(cmdArbiter_io_deqVld),
    .io_deqReady(cmdArbiter_io_deqReady),
    .io_empty(cmdArbiter_io_empty),
    .io_tag(cmdArbiter_io_tag)
  );
  FIFOCore cmdFifos_0 (
    .clock(cmdFifos_0_clock),
    .reset(cmdFifos_0_reset),
    .io_enq_0_addr(cmdFifos_0_io_enq_0_addr),
    .io_enq_0_isWr(cmdFifos_0_io_enq_0_isWr),
    .io_enq_0_size(cmdFifos_0_io_enq_0_size),
    .io_enqVld(cmdFifos_0_io_enqVld),
    .io_deq_0_addr(cmdFifos_0_io_deq_0_addr),
    .io_deq_0_isWr(cmdFifos_0_io_deq_0_isWr),
    .io_deq_0_size(cmdFifos_0_io_deq_0_size),
    .io_deqVld(cmdFifos_0_io_deqVld),
    .io_full(cmdFifos_0_io_full),
    .io_empty(cmdFifos_0_io_empty),
    .io_almostEmpty(cmdFifos_0_io_almostEmpty)
  );
  FIFOCore cmdFifos_1 (
    .clock(cmdFifos_1_clock),
    .reset(cmdFifos_1_reset),
    .io_enq_0_addr(cmdFifos_1_io_enq_0_addr),
    .io_enq_0_isWr(cmdFifos_1_io_enq_0_isWr),
    .io_enq_0_size(cmdFifos_1_io_enq_0_size),
    .io_enqVld(cmdFifos_1_io_enqVld),
    .io_deq_0_addr(cmdFifos_1_io_deq_0_addr),
    .io_deq_0_isWr(cmdFifos_1_io_deq_0_isWr),
    .io_deq_0_size(cmdFifos_1_io_deq_0_size),
    .io_deqVld(cmdFifos_1_io_deqVld),
    .io_full(cmdFifos_1_io_full),
    .io_empty(cmdFifos_1_io_empty),
    .io_almostEmpty(cmdFifos_1_io_almostEmpty)
  );
  FF_136 FF (
    .clock(FF_clock),
    .reset(FF_reset),
    .io_in(FF_io_in),
    .io_init(FF_io_init),
    .io_reset(FF_io_reset),
    .io_out(FF_io_out),
    .io_enable(FF_io_enable)
  );
  Counter_15 sizeCounter (
    .clock(sizeCounter_clock),
    .reset(sizeCounter_reset),
    .io_max(sizeCounter_io_max),
    .io_stride(sizeCounter_io_stride),
    .io_out(sizeCounter_io_out),
    .io_last(sizeCounter_io_last),
    .io_reset(sizeCounter_io_reset),
    .io_enable(sizeCounter_io_enable),
    .io_done(sizeCounter_io_done)
  );
  MuxN_4 isSparseMux (
    .io_ins_0(isSparseMux_io_ins_0),
    .io_ins_1(isSparseMux_io_ins_1),
    .io_sel(isSparseMux_io_sel),
    .io_out(isSparseMux_io_out)
  );
  Counter_15 burstCounter (
    .clock(burstCounter_clock),
    .reset(burstCounter_reset),
    .io_max(burstCounter_io_max),
    .io_stride(burstCounter_io_stride),
    .io_out(burstCounter_io_out),
    .io_last(burstCounter_io_last),
    .io_reset(burstCounter_io_reset),
    .io_enable(burstCounter_io_enable),
    .io_done(burstCounter_io_done)
  );
  Counter_17 burstTagCounter (
    .clock(burstTagCounter_clock),
    .reset(burstTagCounter_reset),
    .io_out(burstTagCounter_io_out),
    .io_reset(burstTagCounter_io_reset),
    .io_enable(burstTagCounter_io_enable)
  );
  FF_115 cmdCooldown (
    .clock(cmdCooldown_clock),
    .reset(cmdCooldown_reset),
    .io_in(cmdCooldown_io_in),
    .io_init(cmdCooldown_io_init),
    .io_reset(cmdCooldown_io_reset),
    .io_out(cmdCooldown_io_out),
    .io_enable(cmdCooldown_io_enable)
  );
  FF_115 burstCounterDoneLatch (
    .clock(burstCounterDoneLatch_clock),
    .reset(burstCounterDoneLatch_reset),
    .io_in(burstCounterDoneLatch_io_in),
    .io_init(burstCounterDoneLatch_io_init),
    .io_reset(burstCounterDoneLatch_io_reset),
    .io_out(burstCounterDoneLatch_io_out),
    .io_enable(burstCounterDoneLatch_io_enable)
  );
  FF_115 sizeCounterDoneLatch (
    .clock(sizeCounterDoneLatch_clock),
    .reset(sizeCounterDoneLatch_reset),
    .io_in(sizeCounterDoneLatch_io_in),
    .io_init(sizeCounterDoneLatch_io_init),
    .io_reset(sizeCounterDoneLatch_io_reset),
    .io_out(sizeCounterDoneLatch_io_out),
    .io_enable(sizeCounterDoneLatch_io_enable)
  );
  MuxN_5 rrespReadyMux (
    .io_ins_0(rrespReadyMux_io_ins_0),
    .io_out(rrespReadyMux_io_out)
  );
  MuxN_6 wdataMux (
    .io_ins_0_valid(wdataMux_io_ins_0_valid),
    .io_ins_0_bits_wdata_0(wdataMux_io_ins_0_bits_wdata_0),
    .io_ins_0_bits_wdata_1(wdataMux_io_ins_0_bits_wdata_1),
    .io_ins_0_bits_wdata_2(wdataMux_io_ins_0_bits_wdata_2),
    .io_ins_0_bits_wdata_3(wdataMux_io_ins_0_bits_wdata_3),
    .io_ins_0_bits_wdata_4(wdataMux_io_ins_0_bits_wdata_4),
    .io_ins_0_bits_wdata_5(wdataMux_io_ins_0_bits_wdata_5),
    .io_ins_0_bits_wdata_6(wdataMux_io_ins_0_bits_wdata_6),
    .io_ins_0_bits_wdata_7(wdataMux_io_ins_0_bits_wdata_7),
    .io_ins_0_bits_wdata_8(wdataMux_io_ins_0_bits_wdata_8),
    .io_ins_0_bits_wdata_9(wdataMux_io_ins_0_bits_wdata_9),
    .io_ins_0_bits_wdata_10(wdataMux_io_ins_0_bits_wdata_10),
    .io_ins_0_bits_wdata_11(wdataMux_io_ins_0_bits_wdata_11),
    .io_ins_0_bits_wdata_12(wdataMux_io_ins_0_bits_wdata_12),
    .io_ins_0_bits_wdata_13(wdataMux_io_ins_0_bits_wdata_13),
    .io_ins_0_bits_wdata_14(wdataMux_io_ins_0_bits_wdata_14),
    .io_ins_0_bits_wdata_15(wdataMux_io_ins_0_bits_wdata_15),
    .io_ins_0_bits_wstrb_0(wdataMux_io_ins_0_bits_wstrb_0),
    .io_ins_0_bits_wstrb_1(wdataMux_io_ins_0_bits_wstrb_1),
    .io_ins_0_bits_wstrb_2(wdataMux_io_ins_0_bits_wstrb_2),
    .io_ins_0_bits_wstrb_3(wdataMux_io_ins_0_bits_wstrb_3),
    .io_ins_0_bits_wstrb_4(wdataMux_io_ins_0_bits_wstrb_4),
    .io_ins_0_bits_wstrb_5(wdataMux_io_ins_0_bits_wstrb_5),
    .io_ins_0_bits_wstrb_6(wdataMux_io_ins_0_bits_wstrb_6),
    .io_ins_0_bits_wstrb_7(wdataMux_io_ins_0_bits_wstrb_7),
    .io_ins_0_bits_wstrb_8(wdataMux_io_ins_0_bits_wstrb_8),
    .io_ins_0_bits_wstrb_9(wdataMux_io_ins_0_bits_wstrb_9),
    .io_ins_0_bits_wstrb_10(wdataMux_io_ins_0_bits_wstrb_10),
    .io_ins_0_bits_wstrb_11(wdataMux_io_ins_0_bits_wstrb_11),
    .io_ins_0_bits_wstrb_12(wdataMux_io_ins_0_bits_wstrb_12),
    .io_ins_0_bits_wstrb_13(wdataMux_io_ins_0_bits_wstrb_13),
    .io_ins_0_bits_wstrb_14(wdataMux_io_ins_0_bits_wstrb_14),
    .io_ins_0_bits_wstrb_15(wdataMux_io_ins_0_bits_wstrb_15),
    .io_ins_0_bits_wstrb_16(wdataMux_io_ins_0_bits_wstrb_16),
    .io_ins_0_bits_wstrb_17(wdataMux_io_ins_0_bits_wstrb_17),
    .io_ins_0_bits_wstrb_18(wdataMux_io_ins_0_bits_wstrb_18),
    .io_ins_0_bits_wstrb_19(wdataMux_io_ins_0_bits_wstrb_19),
    .io_ins_0_bits_wstrb_20(wdataMux_io_ins_0_bits_wstrb_20),
    .io_ins_0_bits_wstrb_21(wdataMux_io_ins_0_bits_wstrb_21),
    .io_ins_0_bits_wstrb_22(wdataMux_io_ins_0_bits_wstrb_22),
    .io_ins_0_bits_wstrb_23(wdataMux_io_ins_0_bits_wstrb_23),
    .io_ins_0_bits_wstrb_24(wdataMux_io_ins_0_bits_wstrb_24),
    .io_ins_0_bits_wstrb_25(wdataMux_io_ins_0_bits_wstrb_25),
    .io_ins_0_bits_wstrb_26(wdataMux_io_ins_0_bits_wstrb_26),
    .io_ins_0_bits_wstrb_27(wdataMux_io_ins_0_bits_wstrb_27),
    .io_ins_0_bits_wstrb_28(wdataMux_io_ins_0_bits_wstrb_28),
    .io_ins_0_bits_wstrb_29(wdataMux_io_ins_0_bits_wstrb_29),
    .io_ins_0_bits_wstrb_30(wdataMux_io_ins_0_bits_wstrb_30),
    .io_ins_0_bits_wstrb_31(wdataMux_io_ins_0_bits_wstrb_31),
    .io_ins_0_bits_wstrb_32(wdataMux_io_ins_0_bits_wstrb_32),
    .io_ins_0_bits_wstrb_33(wdataMux_io_ins_0_bits_wstrb_33),
    .io_ins_0_bits_wstrb_34(wdataMux_io_ins_0_bits_wstrb_34),
    .io_ins_0_bits_wstrb_35(wdataMux_io_ins_0_bits_wstrb_35),
    .io_ins_0_bits_wstrb_36(wdataMux_io_ins_0_bits_wstrb_36),
    .io_ins_0_bits_wstrb_37(wdataMux_io_ins_0_bits_wstrb_37),
    .io_ins_0_bits_wstrb_38(wdataMux_io_ins_0_bits_wstrb_38),
    .io_ins_0_bits_wstrb_39(wdataMux_io_ins_0_bits_wstrb_39),
    .io_ins_0_bits_wstrb_40(wdataMux_io_ins_0_bits_wstrb_40),
    .io_ins_0_bits_wstrb_41(wdataMux_io_ins_0_bits_wstrb_41),
    .io_ins_0_bits_wstrb_42(wdataMux_io_ins_0_bits_wstrb_42),
    .io_ins_0_bits_wstrb_43(wdataMux_io_ins_0_bits_wstrb_43),
    .io_ins_0_bits_wstrb_44(wdataMux_io_ins_0_bits_wstrb_44),
    .io_ins_0_bits_wstrb_45(wdataMux_io_ins_0_bits_wstrb_45),
    .io_ins_0_bits_wstrb_46(wdataMux_io_ins_0_bits_wstrb_46),
    .io_ins_0_bits_wstrb_47(wdataMux_io_ins_0_bits_wstrb_47),
    .io_ins_0_bits_wstrb_48(wdataMux_io_ins_0_bits_wstrb_48),
    .io_ins_0_bits_wstrb_49(wdataMux_io_ins_0_bits_wstrb_49),
    .io_ins_0_bits_wstrb_50(wdataMux_io_ins_0_bits_wstrb_50),
    .io_ins_0_bits_wstrb_51(wdataMux_io_ins_0_bits_wstrb_51),
    .io_ins_0_bits_wstrb_52(wdataMux_io_ins_0_bits_wstrb_52),
    .io_ins_0_bits_wstrb_53(wdataMux_io_ins_0_bits_wstrb_53),
    .io_ins_0_bits_wstrb_54(wdataMux_io_ins_0_bits_wstrb_54),
    .io_ins_0_bits_wstrb_55(wdataMux_io_ins_0_bits_wstrb_55),
    .io_ins_0_bits_wstrb_56(wdataMux_io_ins_0_bits_wstrb_56),
    .io_ins_0_bits_wstrb_57(wdataMux_io_ins_0_bits_wstrb_57),
    .io_ins_0_bits_wstrb_58(wdataMux_io_ins_0_bits_wstrb_58),
    .io_ins_0_bits_wstrb_59(wdataMux_io_ins_0_bits_wstrb_59),
    .io_ins_0_bits_wstrb_60(wdataMux_io_ins_0_bits_wstrb_60),
    .io_ins_0_bits_wstrb_61(wdataMux_io_ins_0_bits_wstrb_61),
    .io_ins_0_bits_wstrb_62(wdataMux_io_ins_0_bits_wstrb_62),
    .io_ins_0_bits_wstrb_63(wdataMux_io_ins_0_bits_wstrb_63),
    .io_out_valid(wdataMux_io_out_valid),
    .io_out_bits_wdata_0(wdataMux_io_out_bits_wdata_0),
    .io_out_bits_wdata_1(wdataMux_io_out_bits_wdata_1),
    .io_out_bits_wdata_2(wdataMux_io_out_bits_wdata_2),
    .io_out_bits_wdata_3(wdataMux_io_out_bits_wdata_3),
    .io_out_bits_wdata_4(wdataMux_io_out_bits_wdata_4),
    .io_out_bits_wdata_5(wdataMux_io_out_bits_wdata_5),
    .io_out_bits_wdata_6(wdataMux_io_out_bits_wdata_6),
    .io_out_bits_wdata_7(wdataMux_io_out_bits_wdata_7),
    .io_out_bits_wdata_8(wdataMux_io_out_bits_wdata_8),
    .io_out_bits_wdata_9(wdataMux_io_out_bits_wdata_9),
    .io_out_bits_wdata_10(wdataMux_io_out_bits_wdata_10),
    .io_out_bits_wdata_11(wdataMux_io_out_bits_wdata_11),
    .io_out_bits_wdata_12(wdataMux_io_out_bits_wdata_12),
    .io_out_bits_wdata_13(wdataMux_io_out_bits_wdata_13),
    .io_out_bits_wdata_14(wdataMux_io_out_bits_wdata_14),
    .io_out_bits_wdata_15(wdataMux_io_out_bits_wdata_15),
    .io_out_bits_wstrb_0(wdataMux_io_out_bits_wstrb_0),
    .io_out_bits_wstrb_1(wdataMux_io_out_bits_wstrb_1),
    .io_out_bits_wstrb_2(wdataMux_io_out_bits_wstrb_2),
    .io_out_bits_wstrb_3(wdataMux_io_out_bits_wstrb_3),
    .io_out_bits_wstrb_4(wdataMux_io_out_bits_wstrb_4),
    .io_out_bits_wstrb_5(wdataMux_io_out_bits_wstrb_5),
    .io_out_bits_wstrb_6(wdataMux_io_out_bits_wstrb_6),
    .io_out_bits_wstrb_7(wdataMux_io_out_bits_wstrb_7),
    .io_out_bits_wstrb_8(wdataMux_io_out_bits_wstrb_8),
    .io_out_bits_wstrb_9(wdataMux_io_out_bits_wstrb_9),
    .io_out_bits_wstrb_10(wdataMux_io_out_bits_wstrb_10),
    .io_out_bits_wstrb_11(wdataMux_io_out_bits_wstrb_11),
    .io_out_bits_wstrb_12(wdataMux_io_out_bits_wstrb_12),
    .io_out_bits_wstrb_13(wdataMux_io_out_bits_wstrb_13),
    .io_out_bits_wstrb_14(wdataMux_io_out_bits_wstrb_14),
    .io_out_bits_wstrb_15(wdataMux_io_out_bits_wstrb_15),
    .io_out_bits_wstrb_16(wdataMux_io_out_bits_wstrb_16),
    .io_out_bits_wstrb_17(wdataMux_io_out_bits_wstrb_17),
    .io_out_bits_wstrb_18(wdataMux_io_out_bits_wstrb_18),
    .io_out_bits_wstrb_19(wdataMux_io_out_bits_wstrb_19),
    .io_out_bits_wstrb_20(wdataMux_io_out_bits_wstrb_20),
    .io_out_bits_wstrb_21(wdataMux_io_out_bits_wstrb_21),
    .io_out_bits_wstrb_22(wdataMux_io_out_bits_wstrb_22),
    .io_out_bits_wstrb_23(wdataMux_io_out_bits_wstrb_23),
    .io_out_bits_wstrb_24(wdataMux_io_out_bits_wstrb_24),
    .io_out_bits_wstrb_25(wdataMux_io_out_bits_wstrb_25),
    .io_out_bits_wstrb_26(wdataMux_io_out_bits_wstrb_26),
    .io_out_bits_wstrb_27(wdataMux_io_out_bits_wstrb_27),
    .io_out_bits_wstrb_28(wdataMux_io_out_bits_wstrb_28),
    .io_out_bits_wstrb_29(wdataMux_io_out_bits_wstrb_29),
    .io_out_bits_wstrb_30(wdataMux_io_out_bits_wstrb_30),
    .io_out_bits_wstrb_31(wdataMux_io_out_bits_wstrb_31),
    .io_out_bits_wstrb_32(wdataMux_io_out_bits_wstrb_32),
    .io_out_bits_wstrb_33(wdataMux_io_out_bits_wstrb_33),
    .io_out_bits_wstrb_34(wdataMux_io_out_bits_wstrb_34),
    .io_out_bits_wstrb_35(wdataMux_io_out_bits_wstrb_35),
    .io_out_bits_wstrb_36(wdataMux_io_out_bits_wstrb_36),
    .io_out_bits_wstrb_37(wdataMux_io_out_bits_wstrb_37),
    .io_out_bits_wstrb_38(wdataMux_io_out_bits_wstrb_38),
    .io_out_bits_wstrb_39(wdataMux_io_out_bits_wstrb_39),
    .io_out_bits_wstrb_40(wdataMux_io_out_bits_wstrb_40),
    .io_out_bits_wstrb_41(wdataMux_io_out_bits_wstrb_41),
    .io_out_bits_wstrb_42(wdataMux_io_out_bits_wstrb_42),
    .io_out_bits_wstrb_43(wdataMux_io_out_bits_wstrb_43),
    .io_out_bits_wstrb_44(wdataMux_io_out_bits_wstrb_44),
    .io_out_bits_wstrb_45(wdataMux_io_out_bits_wstrb_45),
    .io_out_bits_wstrb_46(wdataMux_io_out_bits_wstrb_46),
    .io_out_bits_wstrb_47(wdataMux_io_out_bits_wstrb_47),
    .io_out_bits_wstrb_48(wdataMux_io_out_bits_wstrb_48),
    .io_out_bits_wstrb_49(wdataMux_io_out_bits_wstrb_49),
    .io_out_bits_wstrb_50(wdataMux_io_out_bits_wstrb_50),
    .io_out_bits_wstrb_51(wdataMux_io_out_bits_wstrb_51),
    .io_out_bits_wstrb_52(wdataMux_io_out_bits_wstrb_52),
    .io_out_bits_wstrb_53(wdataMux_io_out_bits_wstrb_53),
    .io_out_bits_wstrb_54(wdataMux_io_out_bits_wstrb_54),
    .io_out_bits_wstrb_55(wdataMux_io_out_bits_wstrb_55),
    .io_out_bits_wstrb_56(wdataMux_io_out_bits_wstrb_56),
    .io_out_bits_wstrb_57(wdataMux_io_out_bits_wstrb_57),
    .io_out_bits_wstrb_58(wdataMux_io_out_bits_wstrb_58),
    .io_out_bits_wstrb_59(wdataMux_io_out_bits_wstrb_59),
    .io_out_bits_wstrb_60(wdataMux_io_out_bits_wstrb_60),
    .io_out_bits_wstrb_61(wdataMux_io_out_bits_wstrb_61),
    .io_out_bits_wstrb_62(wdataMux_io_out_bits_wstrb_62),
    .io_out_bits_wstrb_63(wdataMux_io_out_bits_wstrb_63)
  );
  MuxN_4 cmdDeqValidMux (
    .io_ins_0(cmdDeqValidMux_io_ins_0),
    .io_ins_1(cmdDeqValidMux_io_ins_1),
    .io_sel(cmdDeqValidMux_io_sel),
    .io_out(cmdDeqValidMux_io_out)
  );
  MuxN_8 dramCmdMux (
    .io_ins_0_valid(dramCmdMux_io_ins_0_valid),
    .io_ins_0_bits_addr(dramCmdMux_io_ins_0_bits_addr),
    .io_ins_0_bits_size(dramCmdMux_io_ins_0_bits_size),
    .io_ins_0_bits_isWr(dramCmdMux_io_ins_0_bits_isWr),
    .io_ins_0_bits_tag_uid(dramCmdMux_io_ins_0_bits_tag_uid),
    .io_ins_0_bits_tag_streamId(dramCmdMux_io_ins_0_bits_tag_streamId),
    .io_ins_1_valid(dramCmdMux_io_ins_1_valid),
    .io_ins_1_bits_addr(dramCmdMux_io_ins_1_bits_addr),
    .io_ins_1_bits_size(dramCmdMux_io_ins_1_bits_size),
    .io_ins_1_bits_isWr(dramCmdMux_io_ins_1_bits_isWr),
    .io_ins_1_bits_tag_uid(dramCmdMux_io_ins_1_bits_tag_uid),
    .io_ins_1_bits_tag_streamId(dramCmdMux_io_ins_1_bits_tag_streamId),
    .io_sel(dramCmdMux_io_sel),
    .io_out_valid(dramCmdMux_io_out_valid),
    .io_out_bits_addr(dramCmdMux_io_out_bits_addr),
    .io_out_bits_size(dramCmdMux_io_out_bits_size),
    .io_out_bits_isWr(dramCmdMux_io_out_bits_isWr),
    .io_out_bits_tag_uid(dramCmdMux_io_out_bits_tag_uid),
    .io_out_bits_tag_streamId(dramCmdMux_io_out_bits_tag_streamId)
  );
  FF_143 FF_1 (
    .clock(FF_1_clock),
    .reset(FF_1_reset),
    .io_in(FF_1_io_in),
    .io_out(FF_1_io_out),
    .io_enable(FF_1_io_enable)
  );
  FF_136 FF_2 (
    .clock(FF_2_clock),
    .reset(FF_2_reset),
    .io_in(FF_2_io_in),
    .io_init(FF_2_io_init),
    .io_reset(FF_2_io_reset),
    .io_out(FF_2_io_out),
    .io_enable(FF_2_io_enable)
  );
  FF_145 FF_3 (
    .clock(FF_3_clock),
    .reset(FF_3_reset),
    .io_in(FF_3_io_in),
    .io_out(FF_3_io_out),
    .io_enable(FF_3_io_enable)
  );
  FF_115 FF_4 (
    .clock(FF_4_clock),
    .reset(FF_4_reset),
    .io_in(FF_4_io_in),
    .io_init(FF_4_io_init),
    .io_reset(FF_4_io_reset),
    .io_out(FF_4_io_out),
    .io_enable(FF_4_io_enable)
  );
  FF_137 FF_5 (
    .clock(FF_5_clock),
    .reset(FF_5_reset),
    .io_in(FF_5_io_in),
    .io_out(FF_5_io_out),
    .io_enable(FF_5_io_enable)
  );
  MuxN_5 wrespReadyMux (
    .io_ins_0(wrespReadyMux_io_ins_0),
    .io_out(wrespReadyMux_io_out)
  );
  MuxN_4 gatherLoadIssueMux (
    .io_ins_0(gatherLoadIssueMux_io_ins_0),
    .io_ins_1(gatherLoadIssueMux_io_ins_1),
    .io_sel(gatherLoadIssueMux_io_sel),
    .io_out(gatherLoadIssueMux_io_out)
  );
  Counter_18 gatherLoadIssue (
    .clock(gatherLoadIssue_clock),
    .reset(gatherLoadIssue_reset),
    .io_out(gatherLoadIssue_io_out),
    .io_reset(gatherLoadIssue_io_reset),
    .io_enable(gatherLoadIssue_io_enable)
  );
  MuxN_4 gatherLoadSkipMux (
    .io_ins_0(gatherLoadSkipMux_io_ins_0),
    .io_ins_1(gatherLoadSkipMux_io_ins_1),
    .io_sel(gatherLoadSkipMux_io_sel),
    .io_out(gatherLoadSkipMux_io_out)
  );
  Counter_18 gatherLoadSkip (
    .clock(gatherLoadSkip_clock),
    .reset(gatherLoadSkip_reset),
    .io_out(gatherLoadSkip_io_out),
    .io_reset(gatherLoadSkip_io_reset),
    .io_enable(gatherLoadSkip_io_enable)
  );
  MuxN_4 scatterLoadIssueMux (
    .io_ins_0(scatterLoadIssueMux_io_ins_0),
    .io_ins_1(scatterLoadIssueMux_io_ins_1),
    .io_sel(scatterLoadIssueMux_io_sel),
    .io_out(scatterLoadIssueMux_io_out)
  );
  Counter_18 scatterLoadIssue (
    .clock(scatterLoadIssue_clock),
    .reset(scatterLoadIssue_reset),
    .io_out(scatterLoadIssue_io_out),
    .io_reset(scatterLoadIssue_io_reset),
    .io_enable(scatterLoadIssue_io_enable)
  );
  MuxN_4 scatterLoadSkipMux (
    .io_ins_0(scatterLoadSkipMux_io_ins_0),
    .io_ins_1(scatterLoadSkipMux_io_ins_1),
    .io_sel(scatterLoadSkipMux_io_sel),
    .io_out(scatterLoadSkipMux_io_out)
  );
  Counter_18 scatterLoadSkip (
    .clock(scatterLoadSkip_clock),
    .reset(scatterLoadSkip_reset),
    .io_out(scatterLoadSkip_io_out),
    .io_reset(scatterLoadSkip_io_reset),
    .io_enable(scatterLoadSkip_io_enable)
  );
  MuxN_4 scatterStoreIssueMux (
    .io_ins_0(scatterStoreIssueMux_io_ins_0),
    .io_ins_1(scatterStoreIssueMux_io_ins_1),
    .io_sel(scatterStoreIssueMux_io_sel),
    .io_out(scatterStoreIssueMux_io_out)
  );
  Counter_18 scatterStoreIssue (
    .clock(scatterStoreIssue_clock),
    .reset(scatterStoreIssue_reset),
    .io_out(scatterStoreIssue_io_out),
    .io_reset(scatterStoreIssue_io_reset),
    .io_enable(scatterStoreIssue_io_enable)
  );
  MuxN_4 scatterStoreSkipMux (
    .io_ins_0(scatterStoreSkipMux_io_ins_0),
    .io_ins_1(scatterStoreSkipMux_io_ins_1),
    .io_sel(scatterStoreSkipMux_io_sel),
    .io_out(scatterStoreSkipMux_io_out)
  );
  Counter_18 scatterStoreSkip (
    .clock(scatterStoreSkip_clock),
    .reset(scatterStoreSkip_reset),
    .io_out(scatterStoreSkip_io_out),
    .io_reset(scatterStoreSkip_io_reset),
    .io_enable(scatterStoreSkip_io_enable)
  );
  FIFOWidthConvert denseLoadBuffers_0 (
    .clock(denseLoadBuffers_0_clock),
    .reset(denseLoadBuffers_0_reset),
    .io_enq_0(denseLoadBuffers_0_io_enq_0),
    .io_enq_1(denseLoadBuffers_0_io_enq_1),
    .io_enq_2(denseLoadBuffers_0_io_enq_2),
    .io_enq_3(denseLoadBuffers_0_io_enq_3),
    .io_enq_4(denseLoadBuffers_0_io_enq_4),
    .io_enq_5(denseLoadBuffers_0_io_enq_5),
    .io_enq_6(denseLoadBuffers_0_io_enq_6),
    .io_enq_7(denseLoadBuffers_0_io_enq_7),
    .io_enq_8(denseLoadBuffers_0_io_enq_8),
    .io_enq_9(denseLoadBuffers_0_io_enq_9),
    .io_enq_10(denseLoadBuffers_0_io_enq_10),
    .io_enq_11(denseLoadBuffers_0_io_enq_11),
    .io_enq_12(denseLoadBuffers_0_io_enq_12),
    .io_enq_13(denseLoadBuffers_0_io_enq_13),
    .io_enq_14(denseLoadBuffers_0_io_enq_14),
    .io_enq_15(denseLoadBuffers_0_io_enq_15),
    .io_enqVld(denseLoadBuffers_0_io_enqVld),
    .io_deq_0(denseLoadBuffers_0_io_deq_0),
    .io_deqVld(denseLoadBuffers_0_io_deqVld),
    .io_full(denseLoadBuffers_0_io_full),
    .io_empty(denseLoadBuffers_0_io_empty),
    .io_almostEmpty(denseLoadBuffers_0_io_almostEmpty),
    .io_almostFull(denseLoadBuffers_0_io_almostFull)
  );
  Counter_18 Counter (
    .clock(Counter_clock),
    .reset(Counter_reset),
    .io_out(Counter_io_out),
    .io_reset(Counter_io_reset),
    .io_enable(Counter_io_enable)
  );
  Counter_18 Counter_1 (
    .clock(Counter_1_clock),
    .reset(Counter_1_reset),
    .io_out(Counter_1_io_out),
    .io_reset(Counter_1_io_reset),
    .io_enable(Counter_1_io_enable)
  );
  Counter_18 Counter_2 (
    .clock(Counter_2_clock),
    .reset(Counter_2_reset),
    .io_out(Counter_2_io_out),
    .io_reset(Counter_2_io_reset),
    .io_enable(Counter_2_io_enable)
  );
  Counter_18 Counter_3 (
    .clock(Counter_3_clock),
    .reset(Counter_3_reset),
    .io_out(Counter_3_io_out),
    .io_reset(Counter_3_io_reset),
    .io_enable(Counter_3_io_enable)
  );
  Counter_18 Counter_4 (
    .clock(Counter_4_clock),
    .reset(Counter_4_reset),
    .io_out(Counter_4_io_out),
    .io_reset(Counter_4_io_reset),
    .io_enable(Counter_4_io_enable)
  );
  SRFF SRFF (
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output_data(SRFF_io_output_data)
  );
  SRFF SRFF_1 (
    .clock(SRFF_1_clock),
    .reset(SRFF_1_reset),
    .io_input_set(SRFF_1_io_input_set),
    .io_input_reset(SRFF_1_io_input_reset),
    .io_input_asyn_reset(SRFF_1_io_input_asyn_reset),
    .io_output_data(SRFF_1_io_output_data)
  );
  FF_145 FF_6 (
    .clock(FF_6_clock),
    .reset(FF_6_reset),
    .io_in(FF_6_io_in),
    .io_out(FF_6_io_out),
    .io_enable(FF_6_io_enable)
  );
  FF_180 FF_7 (
    .clock(FF_7_clock),
    .reset(FF_7_reset),
    .io_in(FF_7_io_in),
    .io_out(FF_7_io_out),
    .io_enable(FF_7_io_enable)
  );
  FIFOWidthConvert_1 denseStoreBuffers_0 (
    .clock(denseStoreBuffers_0_clock),
    .reset(denseStoreBuffers_0_reset),
    .io_enqVld(denseStoreBuffers_0_io_enqVld),
    .io_deq_0(denseStoreBuffers_0_io_deq_0),
    .io_deq_1(denseStoreBuffers_0_io_deq_1),
    .io_deq_2(denseStoreBuffers_0_io_deq_2),
    .io_deq_3(denseStoreBuffers_0_io_deq_3),
    .io_deq_4(denseStoreBuffers_0_io_deq_4),
    .io_deq_5(denseStoreBuffers_0_io_deq_5),
    .io_deq_6(denseStoreBuffers_0_io_deq_6),
    .io_deq_7(denseStoreBuffers_0_io_deq_7),
    .io_deq_8(denseStoreBuffers_0_io_deq_8),
    .io_deq_9(denseStoreBuffers_0_io_deq_9),
    .io_deq_10(denseStoreBuffers_0_io_deq_10),
    .io_deq_11(denseStoreBuffers_0_io_deq_11),
    .io_deq_12(denseStoreBuffers_0_io_deq_12),
    .io_deq_13(denseStoreBuffers_0_io_deq_13),
    .io_deq_14(denseStoreBuffers_0_io_deq_14),
    .io_deq_15(denseStoreBuffers_0_io_deq_15),
    .io_deqStrb(denseStoreBuffers_0_io_deqStrb),
    .io_deqVld(denseStoreBuffers_0_io_deqVld),
    .io_full(denseStoreBuffers_0_io_full),
    .io_empty(denseStoreBuffers_0_io_empty),
    .io_almostEmpty(denseStoreBuffers_0_io_almostEmpty),
    .io_almostFull(denseStoreBuffers_0_io_almostFull)
  );
  Counter_15 Counter_5 (
    .clock(Counter_5_clock),
    .reset(Counter_5_reset),
    .io_max(Counter_5_io_max),
    .io_stride(Counter_5_io_stride),
    .io_out(Counter_5_io_out),
    .io_last(Counter_5_io_last),
    .io_reset(Counter_5_io_reset),
    .io_enable(Counter_5_io_enable),
    .io_done(Counter_5_io_done)
  );
  FF_137 FF_8 (
    .clock(FF_8_clock),
    .reset(FF_8_reset),
    .io_in(FF_8_io_in),
    .io_out(FF_8_io_out),
    .io_enable(FF_8_io_enable)
  );
  FIFOCounter FIFOCounter (
    .clock(FIFOCounter_clock),
    .reset(FIFOCounter_reset),
    .io_enqVld(FIFOCounter_io_enqVld),
    .io_full(FIFOCounter_io_full),
    .io_empty(FIFOCounter_io_empty)
  );
  Counter_18 Counter_6 (
    .clock(Counter_6_clock),
    .reset(Counter_6_reset),
    .io_out(Counter_6_io_out),
    .io_reset(Counter_6_io_reset),
    .io_enable(Counter_6_io_enable)
  );
  Counter_18 Counter_7 (
    .clock(Counter_7_clock),
    .reset(Counter_7_reset),
    .io_out(Counter_7_io_out),
    .io_reset(Counter_7_io_reset),
    .io_enable(Counter_7_io_enable)
  );
  Counter_18 Counter_8 (
    .clock(Counter_8_clock),
    .reset(Counter_8_reset),
    .io_out(Counter_8_io_out),
    .io_reset(Counter_8_io_reset),
    .io_enable(Counter_8_io_enable)
  );
  FF_145 burstCounterMaxLatch (
    .clock(burstCounterMaxLatch_clock),
    .reset(burstCounterMaxLatch_reset),
    .io_in(burstCounterMaxLatch_io_in),
    .io_out(burstCounterMaxLatch_io_out),
    .io_enable(burstCounterMaxLatch_io_enable)
  );
  FF_115 dramReadyFF (
    .clock(dramReadyFF_clock),
    .reset(dramReadyFF_reset),
    .io_in(dramReadyFF_io_in),
    .io_init(dramReadyFF_io_init),
    .io_reset(dramReadyFF_io_reset),
    .io_out(dramReadyFF_io_out),
    .io_enable(dramReadyFF_io_enable)
  );
  Counter_18 cycleCount (
    .clock(cycleCount_clock),
    .reset(cycleCount_reset),
    .io_out(cycleCount_io_out),
    .io_reset(cycleCount_io_reset),
    .io_enable(cycleCount_io_enable)
  );
  Counter_18 rdataEnqCount (
    .clock(rdataEnqCount_clock),
    .reset(rdataEnqCount_reset),
    .io_out(rdataEnqCount_io_out),
    .io_reset(rdataEnqCount_io_reset),
    .io_enable(rdataEnqCount_io_enable)
  );
  Counter_18 wdataCount (
    .clock(wdataCount_clock),
    .reset(wdataCount_reset),
    .io_out(wdataCount_io_out),
    .io_reset(wdataCount_io_reset),
    .io_enable(wdataCount_io_enable)
  );
  Counter_18 Counter_9 (
    .clock(Counter_9_clock),
    .reset(Counter_9_reset),
    .io_out(Counter_9_io_out),
    .io_reset(Counter_9_io_reset),
    .io_enable(Counter_9_io_enable)
  );
  Counter_18 Counter_10 (
    .clock(Counter_10_clock),
    .reset(Counter_10_reset),
    .io_out(Counter_10_io_out),
    .io_reset(Counter_10_io_reset),
    .io_enable(Counter_10_io_enable)
  );
  Counter_18 Counter_11 (
    .clock(Counter_11_clock),
    .reset(Counter_11_reset),
    .io_out(Counter_11_io_out),
    .io_reset(Counter_11_io_reset),
    .io_enable(Counter_11_io_enable)
  );
  Counter_18 Counter_12 (
    .clock(Counter_12_clock),
    .reset(Counter_12_reset),
    .io_out(Counter_12_io_out),
    .io_reset(Counter_12_io_reset),
    .io_enable(Counter_12_io_enable)
  );
  Counter_18 Counter_13 (
    .clock(Counter_13_clock),
    .reset(Counter_13_reset),
    .io_out(Counter_13_io_out),
    .io_reset(Counter_13_io_reset),
    .io_enable(Counter_13_io_enable)
  );
  Counter_18 Counter_14 (
    .clock(Counter_14_clock),
    .reset(Counter_14_reset),
    .io_out(Counter_14_io_out),
    .io_reset(Counter_14_io_reset),
    .io_enable(Counter_14_io_enable)
  );
  Counter_18 Counter_15 (
    .clock(Counter_15_clock),
    .reset(Counter_15_reset),
    .io_out(Counter_15_io_out),
    .io_reset(Counter_15_io_reset),
    .io_enable(Counter_15_io_enable)
  );
  Counter_18 Counter_16 (
    .clock(Counter_16_clock),
    .reset(Counter_16_reset),
    .io_out(Counter_16_io_out),
    .io_reset(Counter_16_io_reset),
    .io_enable(Counter_16_io_enable)
  );
  Counter_18 Counter_17 (
    .clock(Counter_17_clock),
    .reset(Counter_17_reset),
    .io_out(Counter_17_io_out),
    .io_reset(Counter_17_io_reset),
    .io_enable(Counter_17_io_enable)
  );
  Counter_18 Counter_18 (
    .clock(Counter_18_clock),
    .reset(Counter_18_reset),
    .io_out(Counter_18_io_out),
    .io_reset(Counter_18_io_reset),
    .io_enable(Counter_18_io_enable)
  );
  Counter_18 Counter_19 (
    .clock(Counter_19_clock),
    .reset(Counter_19_reset),
    .io_out(Counter_19_io_out),
    .io_reset(Counter_19_io_reset),
    .io_enable(Counter_19_io_enable)
  );
  Counter_18 Counter_20 (
    .clock(Counter_20_clock),
    .reset(Counter_20_reset),
    .io_out(Counter_20_io_out),
    .io_reset(Counter_20_io_reset),
    .io_enable(Counter_20_io_enable)
  );
  Counter_18 Counter_21 (
    .clock(Counter_21_clock),
    .reset(Counter_21_reset),
    .io_out(Counter_21_io_out),
    .io_reset(Counter_21_io_reset),
    .io_enable(Counter_21_io_enable)
  );
  Counter_18 Counter_22 (
    .clock(Counter_22_clock),
    .reset(Counter_22_reset),
    .io_out(Counter_22_io_out),
    .io_reset(Counter_22_io_reset),
    .io_enable(Counter_22_io_enable)
  );
  Counter_18 Counter_23 (
    .clock(Counter_23_clock),
    .reset(Counter_23_reset),
    .io_out(Counter_23_io_out),
    .io_reset(Counter_23_io_reset),
    .io_enable(Counter_23_io_enable)
  );
  Counter_18 Counter_24 (
    .clock(Counter_24_clock),
    .reset(Counter_24_reset),
    .io_out(Counter_24_io_out),
    .io_reset(Counter_24_io_reset),
    .io_enable(Counter_24_io_enable)
  );
  Counter_18 Counter_25 (
    .clock(Counter_25_clock),
    .reset(Counter_25_reset),
    .io_out(Counter_25_io_out),
    .io_reset(Counter_25_io_reset),
    .io_enable(Counter_25_io_enable)
  );
  Counter_18 Counter_26 (
    .clock(Counter_26_clock),
    .reset(Counter_26_reset),
    .io_out(Counter_26_io_out),
    .io_reset(Counter_26_io_reset),
    .io_enable(Counter_26_io_enable)
  );
  Counter_18 Counter_27 (
    .clock(Counter_27_clock),
    .reset(Counter_27_reset),
    .io_out(Counter_27_io_out),
    .io_reset(Counter_27_io_reset),
    .io_enable(Counter_27_io_enable)
  );
  Counter_18 Counter_28 (
    .clock(Counter_28_clock),
    .reset(Counter_28_reset),
    .io_out(Counter_28_io_out),
    .io_reset(Counter_28_io_reset),
    .io_enable(Counter_28_io_enable)
  );
  Counter_18 Counter_29 (
    .clock(Counter_29_clock),
    .reset(Counter_29_reset),
    .io_out(Counter_29_io_out),
    .io_reset(Counter_29_io_reset),
    .io_enable(Counter_29_io_enable)
  );
  Counter_18 Counter_30 (
    .clock(Counter_30_clock),
    .reset(Counter_30_reset),
    .io_out(Counter_30_io_out),
    .io_reset(Counter_30_io_reset),
    .io_enable(Counter_30_io_enable)
  );
  Counter_18 Counter_31 (
    .clock(Counter_31_clock),
    .reset(Counter_31_reset),
    .io_out(Counter_31_io_out),
    .io_reset(Counter_31_io_reset),
    .io_enable(Counter_31_io_enable)
  );
  Counter_18 Counter_32 (
    .clock(Counter_32_clock),
    .reset(Counter_32_reset),
    .io_out(Counter_32_io_out),
    .io_reset(Counter_32_io_reset),
    .io_enable(Counter_32_io_enable)
  );
  Counter_18 Counter_33 (
    .clock(Counter_33_clock),
    .reset(Counter_33_reset),
    .io_out(Counter_33_io_out),
    .io_reset(Counter_33_io_reset),
    .io_enable(Counter_33_io_enable)
  );
  Counter_18 Counter_34 (
    .clock(Counter_34_clock),
    .reset(Counter_34_reset),
    .io_out(Counter_34_io_out),
    .io_reset(Counter_34_io_reset),
    .io_enable(Counter_34_io_enable)
  );
  FF_143 FF_9 (
    .clock(FF_9_clock),
    .reset(FF_9_reset),
    .io_in(FF_9_io_in),
    .io_out(FF_9_io_out),
    .io_enable(FF_9_io_enable)
  );
  Counter_18 Counter_35 (
    .clock(Counter_35_clock),
    .reset(Counter_35_reset),
    .io_out(Counter_35_io_out),
    .io_reset(Counter_35_io_reset),
    .io_enable(Counter_35_io_enable)
  );
  Counter_18 Counter_36 (
    .clock(Counter_36_clock),
    .reset(Counter_36_reset),
    .io_out(Counter_36_io_out),
    .io_reset(Counter_36_io_reset),
    .io_enable(Counter_36_io_enable)
  );
  Counter_18 Counter_37 (
    .clock(Counter_37_clock),
    .reset(Counter_37_reset),
    .io_out(Counter_37_io_out),
    .io_reset(Counter_37_io_reset),
    .io_enable(Counter_37_io_enable)
  );
  Counter_18 Counter_38 (
    .clock(Counter_38_clock),
    .reset(Counter_38_reset),
    .io_out(Counter_38_io_out),
    .io_reset(Counter_38_io_reset),
    .io_enable(Counter_38_io_enable)
  );
  Counter_18 Counter_39 (
    .clock(Counter_39_clock),
    .reset(Counter_39_reset),
    .io_out(Counter_39_io_out),
    .io_reset(Counter_39_io_reset),
    .io_enable(Counter_39_io_enable)
  );
  Counter_18 Counter_40 (
    .clock(Counter_40_clock),
    .reset(Counter_40_reset),
    .io_out(Counter_40_io_out),
    .io_reset(Counter_40_io_reset),
    .io_enable(Counter_40_io_enable)
  );
  Counter_18 Counter_41 (
    .clock(Counter_41_clock),
    .reset(Counter_41_reset),
    .io_out(Counter_41_io_out),
    .io_reset(Counter_41_io_reset),
    .io_enable(Counter_41_io_enable)
  );
  Counter_18 Counter_42 (
    .clock(Counter_42_clock),
    .reset(Counter_42_reset),
    .io_out(Counter_42_io_out),
    .io_reset(Counter_42_io_reset),
    .io_enable(Counter_42_io_enable)
  );
  Counter_18 Counter_43 (
    .clock(Counter_43_clock),
    .reset(Counter_43_reset),
    .io_out(Counter_43_io_out),
    .io_reset(Counter_43_io_reset),
    .io_enable(Counter_43_io_enable)
  );
  Counter_18 Counter_44 (
    .clock(Counter_44_clock),
    .reset(Counter_44_reset),
    .io_out(Counter_44_io_out),
    .io_reset(Counter_44_io_reset),
    .io_enable(Counter_44_io_enable)
  );
  Counter_18 Counter_45 (
    .clock(Counter_45_clock),
    .reset(Counter_45_reset),
    .io_out(Counter_45_io_out),
    .io_reset(Counter_45_io_reset),
    .io_enable(Counter_45_io_enable)
  );
  Counter_18 Counter_46 (
    .clock(Counter_46_clock),
    .reset(Counter_46_reset),
    .io_out(Counter_46_io_out),
    .io_reset(Counter_46_io_reset),
    .io_enable(Counter_46_io_enable)
  );
  Counter_18 Counter_47 (
    .clock(Counter_47_clock),
    .reset(Counter_47_reset),
    .io_out(Counter_47_io_out),
    .io_reset(Counter_47_io_reset),
    .io_enable(Counter_47_io_enable)
  );
  Counter_18 Counter_48 (
    .clock(Counter_48_clock),
    .reset(Counter_48_reset),
    .io_out(Counter_48_io_out),
    .io_reset(Counter_48_io_reset),
    .io_enable(Counter_48_io_enable)
  );
  Counter_18 Counter_49 (
    .clock(Counter_49_clock),
    .reset(Counter_49_reset),
    .io_out(Counter_49_io_out),
    .io_reset(Counter_49_io_reset),
    .io_enable(Counter_49_io_enable)
  );
  Counter_18 Counter_50 (
    .clock(Counter_50_clock),
    .reset(Counter_50_reset),
    .io_out(Counter_50_io_out),
    .io_reset(Counter_50_io_reset),
    .io_enable(Counter_50_io_enable)
  );
  Counter_18 Counter_51 (
    .clock(Counter_51_clock),
    .reset(Counter_51_reset),
    .io_out(Counter_51_io_out),
    .io_reset(Counter_51_io_reset),
    .io_enable(Counter_51_io_enable)
  );
  Counter_18 Counter_52 (
    .clock(Counter_52_clock),
    .reset(Counter_52_reset),
    .io_out(Counter_52_io_out),
    .io_reset(Counter_52_io_reset),
    .io_enable(Counter_52_io_enable)
  );
  Counter_18 Counter_53 (
    .clock(Counter_53_clock),
    .reset(Counter_53_reset),
    .io_out(Counter_53_io_out),
    .io_reset(Counter_53_io_reset),
    .io_enable(Counter_53_io_enable)
  );
  Counter_18 Counter_54 (
    .clock(Counter_54_clock),
    .reset(Counter_54_reset),
    .io_out(Counter_54_io_out),
    .io_reset(Counter_54_io_reset),
    .io_enable(Counter_54_io_enable)
  );
  Counter_18 Counter_55 (
    .clock(Counter_55_clock),
    .reset(Counter_55_reset),
    .io_out(Counter_55_io_out),
    .io_reset(Counter_55_io_reset),
    .io_enable(Counter_55_io_enable)
  );
  Counter_18 Counter_56 (
    .clock(Counter_56_clock),
    .reset(Counter_56_reset),
    .io_out(Counter_56_io_out),
    .io_reset(Counter_56_io_reset),
    .io_enable(Counter_56_io_enable)
  );
  Counter_18 Counter_57 (
    .clock(Counter_57_clock),
    .reset(Counter_57_reset),
    .io_out(Counter_57_io_out),
    .io_reset(Counter_57_io_reset),
    .io_enable(Counter_57_io_enable)
  );
  Counter_18 Counter_58 (
    .clock(Counter_58_clock),
    .reset(Counter_58_reset),
    .io_out(Counter_58_io_out),
    .io_reset(Counter_58_io_reset),
    .io_enable(Counter_58_io_enable)
  );
  Counter_18 Counter_59 (
    .clock(Counter_59_clock),
    .reset(Counter_59_reset),
    .io_out(Counter_59_io_out),
    .io_reset(Counter_59_io_reset),
    .io_enable(Counter_59_io_enable)
  );
  FF_136 FF_10 (
    .clock(FF_10_clock),
    .reset(FF_10_reset),
    .io_in(FF_10_io_in),
    .io_init(FF_10_io_init),
    .io_reset(FF_10_io_reset),
    .io_out(FF_10_io_out),
    .io_enable(FF_10_io_enable)
  );
  FF_265 FF_11 (
    .clock(FF_11_clock),
    .reset(FF_11_reset),
    .io_in(FF_11_io_in),
    .io_out(FF_11_io_out),
    .io_enable(FF_11_io_enable)
  );
  FF_266 FF_12 (
    .clock(FF_12_clock),
    .reset(FF_12_reset),
    .io_in(FF_12_io_in),
    .io_out(FF_12_io_out),
    .io_enable(FF_12_io_enable)
  );
  FF_115 FF_13 (
    .clock(FF_13_clock),
    .reset(FF_13_reset),
    .io_in(FF_13_io_in),
    .io_init(FF_13_io_init),
    .io_reset(FF_13_io_reset),
    .io_out(FF_13_io_out),
    .io_enable(FF_13_io_enable)
  );
  FF_268 FF_14 (
    .clock(FF_14_clock),
    .reset(FF_14_reset),
    .io_in(FF_14_io_in),
    .io_out(FF_14_io_out),
    .io_enable(FF_14_io_enable)
  );
  FF_136 FF_15 (
    .clock(FF_15_clock),
    .reset(FF_15_reset),
    .io_in(FF_15_io_in),
    .io_init(FF_15_io_init),
    .io_reset(FF_15_io_reset),
    .io_out(FF_15_io_out),
    .io_enable(FF_15_io_enable)
  );
  FF_265 FF_16 (
    .clock(FF_16_clock),
    .reset(FF_16_reset),
    .io_in(FF_16_io_in),
    .io_out(FF_16_io_out),
    .io_enable(FF_16_io_enable)
  );
  FF_180 FF_17 (
    .clock(FF_17_clock),
    .reset(FF_17_reset),
    .io_in(FF_17_io_in),
    .io_out(FF_17_io_out),
    .io_enable(FF_17_io_enable)
  );
  FF_136 FF_18 (
    .clock(FF_18_clock),
    .reset(FF_18_reset),
    .io_in(FF_18_io_in),
    .io_init(FF_18_io_init),
    .io_reset(FF_18_io_reset),
    .io_out(FF_18_io_out),
    .io_enable(FF_18_io_enable)
  );
  FF_180 FF_19 (
    .clock(FF_19_clock),
    .reset(FF_19_reset),
    .io_in(FF_19_io_in),
    .io_out(FF_19_io_out),
    .io_enable(FF_19_io_enable)
  );
  FF_136 FF_20 (
    .clock(FF_20_clock),
    .reset(FF_20_reset),
    .io_in(FF_20_io_in),
    .io_init(FF_20_io_init),
    .io_reset(FF_20_io_reset),
    .io_out(FF_20_io_out),
    .io_enable(FF_20_io_enable)
  );
  FF_180 FF_21 (
    .clock(FF_21_clock),
    .reset(FF_21_reset),
    .io_in(FF_21_io_in),
    .io_out(FF_21_io_out),
    .io_enable(FF_21_io_enable)
  );
  FF_136 FF_22 (
    .clock(FF_22_clock),
    .reset(FF_22_reset),
    .io_in(FF_22_io_in),
    .io_init(FF_22_io_init),
    .io_reset(FF_22_io_reset),
    .io_out(FF_22_io_out),
    .io_enable(FF_22_io_enable)
  );
  Counter_18 Counter_60 (
    .clock(Counter_60_clock),
    .reset(Counter_60_reset),
    .io_out(Counter_60_io_out),
    .io_reset(Counter_60_io_reset),
    .io_enable(Counter_60_io_enable)
  );
  Counter_18 Counter_61 (
    .clock(Counter_61_clock),
    .reset(Counter_61_reset),
    .io_out(Counter_61_io_out),
    .io_reset(Counter_61_io_reset),
    .io_enable(Counter_61_io_enable)
  );
  Counter_18 Counter_62 (
    .clock(Counter_62_clock),
    .reset(Counter_62_reset),
    .io_out(Counter_62_io_out),
    .io_reset(Counter_62_io_reset),
    .io_enable(Counter_62_io_enable)
  );
  Counter_18 Counter_63 (
    .clock(Counter_63_clock),
    .reset(Counter_63_reset),
    .io_out(Counter_63_io_out),
    .io_reset(Counter_63_io_reset),
    .io_enable(Counter_63_io_enable)
  );
  Counter_18 Counter_64 (
    .clock(Counter_64_clock),
    .reset(Counter_64_reset),
    .io_out(Counter_64_io_out),
    .io_reset(Counter_64_io_reset),
    .io_enable(Counter_64_io_enable)
  );
  Counter_18 Counter_65 (
    .clock(Counter_65_clock),
    .reset(Counter_65_reset),
    .io_out(Counter_65_io_out),
    .io_reset(Counter_65_io_reset),
    .io_enable(Counter_65_io_enable)
  );
  Counter_18 Counter_66 (
    .clock(Counter_66_clock),
    .reset(Counter_66_reset),
    .io_out(Counter_66_io_out),
    .io_reset(Counter_66_io_reset),
    .io_enable(Counter_66_io_enable)
  );
  Counter_18 Counter_67 (
    .clock(Counter_67_clock),
    .reset(Counter_67_reset),
    .io_out(Counter_67_io_out),
    .io_reset(Counter_67_io_reset),
    .io_enable(Counter_67_io_enable)
  );
  Counter_18 Counter_68 (
    .clock(Counter_68_clock),
    .reset(Counter_68_reset),
    .io_out(Counter_68_io_out),
    .io_reset(Counter_68_io_reset),
    .io_enable(Counter_68_io_enable)
  );
  Counter_18 Counter_69 (
    .clock(Counter_69_clock),
    .reset(Counter_69_reset),
    .io_out(Counter_69_io_out),
    .io_reset(Counter_69_io_reset),
    .io_enable(Counter_69_io_enable)
  );
  Counter_18 Counter_70 (
    .clock(Counter_70_clock),
    .reset(Counter_70_reset),
    .io_out(Counter_70_io_out),
    .io_reset(Counter_70_io_reset),
    .io_enable(Counter_70_io_enable)
  );
  Counter_18 Counter_71 (
    .clock(Counter_71_clock),
    .reset(Counter_71_reset),
    .io_out(Counter_71_io_out),
    .io_reset(Counter_71_io_reset),
    .io_enable(Counter_71_io_enable)
  );
  Counter_18 Counter_72 (
    .clock(Counter_72_clock),
    .reset(Counter_72_reset),
    .io_out(Counter_72_io_out),
    .io_reset(Counter_72_io_reset),
    .io_enable(Counter_72_io_enable)
  );
  FF_136 FF_23 (
    .clock(FF_23_clock),
    .reset(FF_23_reset),
    .io_in(FF_23_io_in),
    .io_init(FF_23_io_init),
    .io_reset(FF_23_io_reset),
    .io_out(FF_23_io_out),
    .io_enable(FF_23_io_enable)
  );
  FF_265 FF_24 (
    .clock(FF_24_clock),
    .reset(FF_24_reset),
    .io_in(FF_24_io_in),
    .io_out(FF_24_io_out),
    .io_enable(FF_24_io_enable)
  );
  FF_266 FF_25 (
    .clock(FF_25_clock),
    .reset(FF_25_reset),
    .io_in(FF_25_io_in),
    .io_out(FF_25_io_out),
    .io_enable(FF_25_io_enable)
  );
  FF_268 FF_26 (
    .clock(FF_26_clock),
    .reset(FF_26_reset),
    .io_in(FF_26_io_in),
    .io_out(FF_26_io_out),
    .io_enable(FF_26_io_enable)
  );
  FF_136 FF_27 (
    .clock(FF_27_clock),
    .reset(FF_27_reset),
    .io_in(FF_27_io_in),
    .io_init(FF_27_io_init),
    .io_reset(FF_27_io_reset),
    .io_out(FF_27_io_out),
    .io_enable(FF_27_io_enable)
  );
  FF_265 FF_28 (
    .clock(FF_28_clock),
    .reset(FF_28_reset),
    .io_in(FF_28_io_in),
    .io_out(FF_28_io_out),
    .io_enable(FF_28_io_enable)
  );
  FF_180 FF_29 (
    .clock(FF_29_clock),
    .reset(FF_29_reset),
    .io_in(FF_29_io_in),
    .io_out(FF_29_io_out),
    .io_enable(FF_29_io_enable)
  );
  FF_136 FF_30 (
    .clock(FF_30_clock),
    .reset(FF_30_reset),
    .io_in(FF_30_io_in),
    .io_init(FF_30_io_init),
    .io_reset(FF_30_io_reset),
    .io_out(FF_30_io_out),
    .io_enable(FF_30_io_enable)
  );
  FF_180 FF_31 (
    .clock(FF_31_clock),
    .reset(FF_31_reset),
    .io_in(FF_31_io_in),
    .io_out(FF_31_io_out),
    .io_enable(FF_31_io_enable)
  );
  FF_136 FF_32 (
    .clock(FF_32_clock),
    .reset(FF_32_reset),
    .io_in(FF_32_io_in),
    .io_init(FF_32_io_init),
    .io_reset(FF_32_io_reset),
    .io_out(FF_32_io_out),
    .io_enable(FF_32_io_enable)
  );
  FF_180 FF_33 (
    .clock(FF_33_clock),
    .reset(FF_33_reset),
    .io_in(FF_33_io_in),
    .io_out(FF_33_io_out),
    .io_enable(FF_33_io_enable)
  );
  FF_136 FF_34 (
    .clock(FF_34_clock),
    .reset(FF_34_reset),
    .io_in(FF_34_io_in),
    .io_init(FF_34_io_init),
    .io_reset(FF_34_io_reset),
    .io_out(FF_34_io_out),
    .io_enable(FF_34_io_enable)
  );
  assign _T_886 = io_app_loads_0_cmd_bits_addr[31:0];
  assign _T_887 = {32'h7f,_T_886};
  assign _T_891 = ~ cmdArbiter_io_full_0;
  assign _GEN_0 = {{48'd0}, sizeCounter_io_out};
  assign _T_894 = cmdArbiter_io_deq_0_addr + _GEN_0;
  assign _T_895 = _T_894[63:0];
  assign _T_896 = io_enable & cmdArbiter_io_deqReady;
  assign _T_897 = ~ cmdArbiter_io_deq_0_isWr;
  assign cmdRead = _T_896 & _T_897;
  assign cmdWrite = _T_896 & cmdArbiter_io_deq_0_isWr;
  assign _T_903 = isSparseMux_io_out ? 16'h1 : cmdArbiter_io_deq_0_size;
  assign _T_908 = isSparseMux_io_out ? 1'h0 : sizeCounter_io_done;
  assign _T_931 = cmdAddr_bits[63:6];
  assign _T_933 = {_T_931,6'h0};
  assign _T_938 = cmdArbiter_io_deq_0_size - sizeCounter_io_out;
  assign _T_939 = $unsigned(_T_938);
  assign _T_940 = _T_939[15:0];
  assign _T_942 = sizeCounter_io_done ? _T_940 : 16'h4000;
  assign _T_943 = isSparseMux_io_out ? cmdArbiter_io_deq_0_size : _T_942;
  assign _T_944 = _T_937_bits[15:6];
  assign _T_945 = _T_937_bits[5:0];
  assign _T_947 = _T_945 != 6'h0;
  assign _GEN_2 = {{9'd0}, _T_947};
  assign _T_948 = _T_944 + _GEN_2;
  assign _T_949 = _T_948[9:0];
  assign _T_950 = ~ dramCmdMux_io_out_bits_isWr;
  assign _T_951 = dramCmdMux_io_out_valid & _T_950;
  assign _T_978 = _T_971_bits[15:6];
  assign _T_979 = _T_971_bits[5:0];
  assign _T_981 = _T_979 != 6'h0;
  assign _GEN_3 = {{9'd0}, _T_981};
  assign _T_982 = _T_978 + _GEN_3;
  assign _T_983 = _T_982[9:0];
  assign _T_1027 = io_dram_rresp_bits_tag_streamId == 6'h0;
  assign _T_1028 = io_dram_rresp_valid & _T_1027;
  assign _T_1029 = ~ denseLoadBuffers_0_io_full;
  assign _T_1031 = ~ denseLoadBuffers_0_io_empty;
  assign _T_1046 = _T_1031 & io_app_loads_0_rdata_ready;
  assign _T_1051 = denseLoadBuffers_0_io_empty & denseLoadBuffers_0_io_deqVld;
  assign _T_1057 = reset | io_reset;
  assign _T_1064 = ~ SRFF_io_output_data;
  assign _T_1065 = ~ denseLoadBuffers_0_io_deqVld;
  assign _T_1074 = denseLoadBuffers_0_io_deqVld & _T_1068;
  assign _T_1075 = _T_1064 & _T_1074;
  assign _T_1079 = ~ SRFF_1_io_output_data;
  assign _T_1080 = ~ denseLoadBuffers_0_io_enqVld;
  assign _T_1089 = denseLoadBuffers_0_io_enqVld & _T_1083;
  assign _T_1090 = _T_1079 & _T_1089;
  assign _T_1091 = {denseLoadBuffers_0_io_enq_15,denseLoadBuffers_0_io_enq_14};
  assign _T_1092 = {_T_1091,denseLoadBuffers_0_io_enq_13};
  assign _T_1093 = {_T_1092,denseLoadBuffers_0_io_enq_12};
  assign _T_1094 = {_T_1093,denseLoadBuffers_0_io_enq_11};
  assign _T_1095 = {_T_1094,denseLoadBuffers_0_io_enq_10};
  assign _T_1096 = {_T_1095,denseLoadBuffers_0_io_enq_9};
  assign _T_1097 = {_T_1096,denseLoadBuffers_0_io_enq_8};
  assign _T_1098 = {_T_1097,denseLoadBuffers_0_io_enq_7};
  assign _T_1099 = {_T_1098,denseLoadBuffers_0_io_enq_6};
  assign _T_1100 = {_T_1099,denseLoadBuffers_0_io_enq_5};
  assign _T_1101 = {_T_1100,denseLoadBuffers_0_io_enq_4};
  assign _T_1102 = {_T_1101,denseLoadBuffers_0_io_enq_3};
  assign _T_1103 = {_T_1102,denseLoadBuffers_0_io_enq_2};
  assign _T_1104 = {_T_1103,denseLoadBuffers_0_io_enq_1};
  assign _T_1105 = {_T_1104,denseLoadBuffers_0_io_enq_0};
  assign _T_1109 = burstCounterDoneLatch_io_out & sizeCounterDoneLatch_io_out;
  assign _T_1110 = cmdWrite & wdataMux_io_out_valid;
  assign _T_1111 = ~ dramReadySeen;
  assign _T_1112 = _T_1110 & _T_1111;
  assign _T_1114 = ~ denseStoreBuffers_0_io_empty;
  assign _T_1115 = cmdWrite & _T_1114;
  assign _T_1116 = _T_1115 & io_dram_wdata_ready;
  assign _T_1118 = cmdArbiter_io_tag;
  assign _T_1119 = _T_1116 & _T_1118;
  assign _T_1120 = ~ cmdCooldown_io_out;
  assign _T_1121 = _T_1119 & _T_1120;
  assign _T_1122 = ~ burstCounterDoneLatch_io_out;
  assign _T_1123 = _T_1121 & _T_1122;
  assign _T_1127 = _T_1115 & _T_1120;
  assign _T_1129 = _T_1127 & _T_1122;
  assign _T_1130 = denseStoreBuffers_0_io_deqStrb[0];
  assign _T_1131 = denseStoreBuffers_0_io_deqStrb[1];
  assign _T_1132 = denseStoreBuffers_0_io_deqStrb[2];
  assign _T_1133 = denseStoreBuffers_0_io_deqStrb[3];
  assign _T_1134 = denseStoreBuffers_0_io_deqStrb[4];
  assign _T_1135 = denseStoreBuffers_0_io_deqStrb[5];
  assign _T_1136 = denseStoreBuffers_0_io_deqStrb[6];
  assign _T_1137 = denseStoreBuffers_0_io_deqStrb[7];
  assign _T_1138 = denseStoreBuffers_0_io_deqStrb[8];
  assign _T_1139 = denseStoreBuffers_0_io_deqStrb[9];
  assign _T_1140 = denseStoreBuffers_0_io_deqStrb[10];
  assign _T_1141 = denseStoreBuffers_0_io_deqStrb[11];
  assign _T_1142 = denseStoreBuffers_0_io_deqStrb[12];
  assign _T_1143 = denseStoreBuffers_0_io_deqStrb[13];
  assign _T_1144 = denseStoreBuffers_0_io_deqStrb[14];
  assign _T_1145 = denseStoreBuffers_0_io_deqStrb[15];
  assign _T_1146 = denseStoreBuffers_0_io_deqStrb[16];
  assign _T_1147 = denseStoreBuffers_0_io_deqStrb[17];
  assign _T_1148 = denseStoreBuffers_0_io_deqStrb[18];
  assign _T_1149 = denseStoreBuffers_0_io_deqStrb[19];
  assign _T_1150 = denseStoreBuffers_0_io_deqStrb[20];
  assign _T_1151 = denseStoreBuffers_0_io_deqStrb[21];
  assign _T_1152 = denseStoreBuffers_0_io_deqStrb[22];
  assign _T_1153 = denseStoreBuffers_0_io_deqStrb[23];
  assign _T_1154 = denseStoreBuffers_0_io_deqStrb[24];
  assign _T_1155 = denseStoreBuffers_0_io_deqStrb[25];
  assign _T_1156 = denseStoreBuffers_0_io_deqStrb[26];
  assign _T_1157 = denseStoreBuffers_0_io_deqStrb[27];
  assign _T_1158 = denseStoreBuffers_0_io_deqStrb[28];
  assign _T_1159 = denseStoreBuffers_0_io_deqStrb[29];
  assign _T_1160 = denseStoreBuffers_0_io_deqStrb[30];
  assign _T_1161 = denseStoreBuffers_0_io_deqStrb[31];
  assign _T_1162 = denseStoreBuffers_0_io_deqStrb[32];
  assign _T_1163 = denseStoreBuffers_0_io_deqStrb[33];
  assign _T_1164 = denseStoreBuffers_0_io_deqStrb[34];
  assign _T_1165 = denseStoreBuffers_0_io_deqStrb[35];
  assign _T_1166 = denseStoreBuffers_0_io_deqStrb[36];
  assign _T_1167 = denseStoreBuffers_0_io_deqStrb[37];
  assign _T_1168 = denseStoreBuffers_0_io_deqStrb[38];
  assign _T_1169 = denseStoreBuffers_0_io_deqStrb[39];
  assign _T_1170 = denseStoreBuffers_0_io_deqStrb[40];
  assign _T_1171 = denseStoreBuffers_0_io_deqStrb[41];
  assign _T_1172 = denseStoreBuffers_0_io_deqStrb[42];
  assign _T_1173 = denseStoreBuffers_0_io_deqStrb[43];
  assign _T_1174 = denseStoreBuffers_0_io_deqStrb[44];
  assign _T_1175 = denseStoreBuffers_0_io_deqStrb[45];
  assign _T_1176 = denseStoreBuffers_0_io_deqStrb[46];
  assign _T_1177 = denseStoreBuffers_0_io_deqStrb[47];
  assign _T_1178 = denseStoreBuffers_0_io_deqStrb[48];
  assign _T_1179 = denseStoreBuffers_0_io_deqStrb[49];
  assign _T_1180 = denseStoreBuffers_0_io_deqStrb[50];
  assign _T_1181 = denseStoreBuffers_0_io_deqStrb[51];
  assign _T_1182 = denseStoreBuffers_0_io_deqStrb[52];
  assign _T_1183 = denseStoreBuffers_0_io_deqStrb[53];
  assign _T_1184 = denseStoreBuffers_0_io_deqStrb[54];
  assign _T_1185 = denseStoreBuffers_0_io_deqStrb[55];
  assign _T_1186 = denseStoreBuffers_0_io_deqStrb[56];
  assign _T_1187 = denseStoreBuffers_0_io_deqStrb[57];
  assign _T_1188 = denseStoreBuffers_0_io_deqStrb[58];
  assign _T_1189 = denseStoreBuffers_0_io_deqStrb[59];
  assign _T_1190 = denseStoreBuffers_0_io_deqStrb[60];
  assign _T_1191 = denseStoreBuffers_0_io_deqStrb[61];
  assign _T_1192 = denseStoreBuffers_0_io_deqStrb[62];
  assign _T_1193 = denseStoreBuffers_0_io_deqStrb[63];
  assign _T_1194 = ~ denseStoreBuffers_0_io_full;
  assign _T_1197 = io_dram_cmd_valid & io_dram_cmd_ready;
  assign _T_1202 = io_dram_wresp_bits_tag_streamId == 6'h1;
  assign _T_1203 = io_dram_wresp_valid & _T_1202;
  assign _T_1204 = ~ FIFOCounter_io_full;
  assign _T_1205 = ~ FIFOCounter_io_empty;
  assign burstCounterMax = _T_1197 ? io_dram_cmd_bits_size : burstCounterMaxLatch_io_out;
  assign _T_1227 = isSparseMux_io_out ? 1'h0 : burstCounter_io_done;
  assign _T_1229 = burstCounter_io_last ? _T_1109 : burstCounterDoneLatch_io_out;
  assign _T_1231 = io_dram_cmd_bits_isWr ? burstCounterMax : 32'h1;
  assign _T_1233 = wdataMux_io_out_valid & io_dram_wdata_ready;
  assign _T_1235 = io_dram_cmd_bits_isWr ? _T_1233 : _T_1197;
  assign dramReadyFFEnabler = isSparseMux_io_out ? burstCounter_io_done : burstCounterDoneLatch_io_out;
  assign _T_1243 = io_dram_cmd_valid & io_dram_cmd_bits_isWr;
  assign _T_1244 = dramReadyFFEnabler | _T_1243;
  assign _T_1246 = io_dram_cmd_ready | dramReadySeen;
  assign _T_1247 = dramReadyFFEnabler ? 1'h0 : _T_1246;
  assign _T_1249 = ~ _T_1197;
  assign _T_1255 = isSparseMux_io_out ? 1'h1 : _T_1120;
  assign _T_1256 = dramCmdMux_io_out_valid & _T_1255;
  assign _T_1261 = io_dram_rresp_valid & io_dram_rresp_ready;
  assign _T_1266 = io_dram_wdata_valid & io_dram_wdata_ready;
  assign _T_1267 = _T_1266 & io_enable;
  assign _T_1272 = io_enable & io_dram_cmd_ready;
  assign _T_1273 = _T_1272 & io_dram_cmd_valid;
  assign _T_1278 = ~ cmdArbiter_io_empty;
  assign _T_1279 = io_enable & _T_1278;
  assign _T_1280 = io_dram_cmd_ready & io_dram_cmd_valid;
  assign _T_1281 = ~ _T_1280;
  assign _T_1282 = _T_1279 & _T_1281;
  assign _T_1290 = _T_1273 & _T_897;
  assign _T_1295 = io_enable & io_app_loads_0_cmd_valid;
  assign _T_1301 = _T_1295 & io_app_loads_0_cmd_ready;
  assign _T_1308 = cmdArbiter_io_tag == 1'h0;
  assign _T_1309 = _T_1197 & _T_1308;
  assign _T_1316 = _T_1273 & cmdArbiter_io_deq_0_isWr;
  assign _T_1335 = _T_1197 & _T_1118;
  assign _T_1345 = io_enable & io_dram_rresp_valid;
  assign _T_1346 = ~ io_dram_rresp_ready;
  assign _T_1347 = _T_1345 & _T_1346;
  assign _T_1352 = ~ io_dram_rresp_valid;
  assign _T_1353 = io_enable & _T_1352;
  assign _T_1354 = _T_1353 & io_dram_rresp_ready;
  assign _T_1362 = _T_1261 & _T_1027;
  assign _T_1367 = io_dram_wresp_valid & io_dram_wresp_ready;
  assign _T_1372 = io_enable & io_dram_wresp_valid;
  assign _T_1373 = ~ io_dram_wresp_ready;
  assign _T_1374 = _T_1372 & _T_1373;
  assign _T_1379 = ~ io_dram_wresp_valid;
  assign _T_1380 = io_enable & _T_1379;
  assign _T_1381 = _T_1380 & io_dram_wresp_ready;
  assign _T_1389 = _T_1367 & _T_1202;
  assign _T_1425 = io_dram_rresp_bits_tag_streamId >= 6'h1;
  assign _T_1443 = _T_1194 & denseStoreBuffers_0_io_enqVld;
  assign _T_1448 = denseStoreBuffers_0_io_full & denseStoreBuffers_0_io_enqVld;
  assign _T_1469 = io_dram_rresp_valid & denseLoadBuffers_0_io_enqVld;
  assign _T_1480 = _T_1261 & denseLoadBuffers_0_io_enqVld;
  assign _T_1486 = io_dram_rresp_valid & _T_1346;
  assign _T_1499 = io_TOP_AXI_ARREADY & io_TOP_AXI_ARVALID;
  assign _T_1508 = io_TOP_AXI_AWREADY & io_TOP_AXI_AWVALID;
  assign _T_1517 = io_TOP_AXI_RREADY & io_TOP_AXI_RVALID;
  assign _T_1526 = io_TOP_AXI_WREADY & io_TOP_AXI_WVALID;
  assign _T_1531 = ~ io_TOP_AXI_WREADY;
  assign _T_1532 = _T_1531 & io_TOP_AXI_WVALID;
  assign _T_1546 = io_TOP_AXI_BREADY & io_TOP_AXI_BVALID;
  assign _T_1551 = io_TOP_AXI_ARVALID & io_TOP_AXI_ARREADY;
  assign _T_1571 = io_TOP_AXI_AWVALID & io_TOP_AXI_AWREADY;
  assign _T_1579 = io_TOP_AXI_WVALID & io_TOP_AXI_WREADY;
  assign _T_1589 = wdataCount_io_out == 64'h0;
  assign _T_1590 = _T_1579 & _T_1589;
  assign _T_1603 = wdataCount_io_out == 64'h1;
  assign _T_1604 = _T_1579 & _T_1603;
  assign _T_1623 = io_DWIDTH_AXI_ARREADY & io_DWIDTH_AXI_ARVALID;
  assign _T_1632 = io_DWIDTH_AXI_AWREADY & io_DWIDTH_AXI_AWVALID;
  assign _T_1641 = io_DWIDTH_AXI_RREADY & io_DWIDTH_AXI_RVALID;
  assign _T_1650 = io_DWIDTH_AXI_WREADY & io_DWIDTH_AXI_WVALID;
  assign _T_1655 = ~ io_DWIDTH_AXI_WREADY;
  assign _T_1656 = _T_1655 & io_DWIDTH_AXI_WVALID;
  assign _T_1670 = io_DWIDTH_AXI_BREADY & io_DWIDTH_AXI_BVALID;
  assign _T_1675 = io_DWIDTH_AXI_ARVALID & io_DWIDTH_AXI_ARREADY;
  assign _T_1691 = io_DWIDTH_AXI_AWVALID & io_DWIDTH_AXI_AWREADY;
  assign _T_1699 = io_DWIDTH_AXI_WVALID & io_DWIDTH_AXI_WREADY;
  assign _T_1710 = _T_1699 & _T_1589;
  assign _T_1724 = _T_1699 & _T_1603;
  assign io_app_loads_0_cmd_ready = _T_891;
  assign io_app_loads_0_rdata_valid = _T_1031;
  assign io_app_loads_0_rdata_bits_0 = denseLoadBuffers_0_io_deq_0;
  assign io_dram_cmd_valid = _T_1256;
  assign io_dram_cmd_bits_addr = dramCmdMux_io_out_bits_addr;
  assign io_dram_cmd_bits_size = dramCmdMux_io_out_bits_size;
  assign io_dram_cmd_bits_isWr = dramCmdMux_io_out_bits_isWr;
  assign io_dram_cmd_bits_tag_uid = dramCmdMux_io_out_bits_tag_uid;
  assign io_dram_cmd_bits_tag_streamId = dramCmdMux_io_out_bits_tag_streamId;
  assign io_dram_wdata_valid = wdataMux_io_out_valid;
  assign io_dram_wdata_bits_wdata_0 = wdataMux_io_out_bits_wdata_0;
  assign io_dram_wdata_bits_wdata_1 = wdataMux_io_out_bits_wdata_1;
  assign io_dram_wdata_bits_wdata_2 = wdataMux_io_out_bits_wdata_2;
  assign io_dram_wdata_bits_wdata_3 = wdataMux_io_out_bits_wdata_3;
  assign io_dram_wdata_bits_wdata_4 = wdataMux_io_out_bits_wdata_4;
  assign io_dram_wdata_bits_wdata_5 = wdataMux_io_out_bits_wdata_5;
  assign io_dram_wdata_bits_wdata_6 = wdataMux_io_out_bits_wdata_6;
  assign io_dram_wdata_bits_wdata_7 = wdataMux_io_out_bits_wdata_7;
  assign io_dram_wdata_bits_wdata_8 = wdataMux_io_out_bits_wdata_8;
  assign io_dram_wdata_bits_wdata_9 = wdataMux_io_out_bits_wdata_9;
  assign io_dram_wdata_bits_wdata_10 = wdataMux_io_out_bits_wdata_10;
  assign io_dram_wdata_bits_wdata_11 = wdataMux_io_out_bits_wdata_11;
  assign io_dram_wdata_bits_wdata_12 = wdataMux_io_out_bits_wdata_12;
  assign io_dram_wdata_bits_wdata_13 = wdataMux_io_out_bits_wdata_13;
  assign io_dram_wdata_bits_wdata_14 = wdataMux_io_out_bits_wdata_14;
  assign io_dram_wdata_bits_wdata_15 = wdataMux_io_out_bits_wdata_15;
  assign io_dram_wdata_bits_wstrb_0 = wdataMux_io_out_bits_wstrb_63;
  assign io_dram_wdata_bits_wstrb_1 = wdataMux_io_out_bits_wstrb_62;
  assign io_dram_wdata_bits_wstrb_2 = wdataMux_io_out_bits_wstrb_61;
  assign io_dram_wdata_bits_wstrb_3 = wdataMux_io_out_bits_wstrb_60;
  assign io_dram_wdata_bits_wstrb_4 = wdataMux_io_out_bits_wstrb_59;
  assign io_dram_wdata_bits_wstrb_5 = wdataMux_io_out_bits_wstrb_58;
  assign io_dram_wdata_bits_wstrb_6 = wdataMux_io_out_bits_wstrb_57;
  assign io_dram_wdata_bits_wstrb_7 = wdataMux_io_out_bits_wstrb_56;
  assign io_dram_wdata_bits_wstrb_8 = wdataMux_io_out_bits_wstrb_55;
  assign io_dram_wdata_bits_wstrb_9 = wdataMux_io_out_bits_wstrb_54;
  assign io_dram_wdata_bits_wstrb_10 = wdataMux_io_out_bits_wstrb_53;
  assign io_dram_wdata_bits_wstrb_11 = wdataMux_io_out_bits_wstrb_52;
  assign io_dram_wdata_bits_wstrb_12 = wdataMux_io_out_bits_wstrb_51;
  assign io_dram_wdata_bits_wstrb_13 = wdataMux_io_out_bits_wstrb_50;
  assign io_dram_wdata_bits_wstrb_14 = wdataMux_io_out_bits_wstrb_49;
  assign io_dram_wdata_bits_wstrb_15 = wdataMux_io_out_bits_wstrb_48;
  assign io_dram_wdata_bits_wstrb_16 = wdataMux_io_out_bits_wstrb_47;
  assign io_dram_wdata_bits_wstrb_17 = wdataMux_io_out_bits_wstrb_46;
  assign io_dram_wdata_bits_wstrb_18 = wdataMux_io_out_bits_wstrb_45;
  assign io_dram_wdata_bits_wstrb_19 = wdataMux_io_out_bits_wstrb_44;
  assign io_dram_wdata_bits_wstrb_20 = wdataMux_io_out_bits_wstrb_43;
  assign io_dram_wdata_bits_wstrb_21 = wdataMux_io_out_bits_wstrb_42;
  assign io_dram_wdata_bits_wstrb_22 = wdataMux_io_out_bits_wstrb_41;
  assign io_dram_wdata_bits_wstrb_23 = wdataMux_io_out_bits_wstrb_40;
  assign io_dram_wdata_bits_wstrb_24 = wdataMux_io_out_bits_wstrb_39;
  assign io_dram_wdata_bits_wstrb_25 = wdataMux_io_out_bits_wstrb_38;
  assign io_dram_wdata_bits_wstrb_26 = wdataMux_io_out_bits_wstrb_37;
  assign io_dram_wdata_bits_wstrb_27 = wdataMux_io_out_bits_wstrb_36;
  assign io_dram_wdata_bits_wstrb_28 = wdataMux_io_out_bits_wstrb_35;
  assign io_dram_wdata_bits_wstrb_29 = wdataMux_io_out_bits_wstrb_34;
  assign io_dram_wdata_bits_wstrb_30 = wdataMux_io_out_bits_wstrb_33;
  assign io_dram_wdata_bits_wstrb_31 = wdataMux_io_out_bits_wstrb_32;
  assign io_dram_wdata_bits_wstrb_32 = wdataMux_io_out_bits_wstrb_31;
  assign io_dram_wdata_bits_wstrb_33 = wdataMux_io_out_bits_wstrb_30;
  assign io_dram_wdata_bits_wstrb_34 = wdataMux_io_out_bits_wstrb_29;
  assign io_dram_wdata_bits_wstrb_35 = wdataMux_io_out_bits_wstrb_28;
  assign io_dram_wdata_bits_wstrb_36 = wdataMux_io_out_bits_wstrb_27;
  assign io_dram_wdata_bits_wstrb_37 = wdataMux_io_out_bits_wstrb_26;
  assign io_dram_wdata_bits_wstrb_38 = wdataMux_io_out_bits_wstrb_25;
  assign io_dram_wdata_bits_wstrb_39 = wdataMux_io_out_bits_wstrb_24;
  assign io_dram_wdata_bits_wstrb_40 = wdataMux_io_out_bits_wstrb_23;
  assign io_dram_wdata_bits_wstrb_41 = wdataMux_io_out_bits_wstrb_22;
  assign io_dram_wdata_bits_wstrb_42 = wdataMux_io_out_bits_wstrb_21;
  assign io_dram_wdata_bits_wstrb_43 = wdataMux_io_out_bits_wstrb_20;
  assign io_dram_wdata_bits_wstrb_44 = wdataMux_io_out_bits_wstrb_19;
  assign io_dram_wdata_bits_wstrb_45 = wdataMux_io_out_bits_wstrb_18;
  assign io_dram_wdata_bits_wstrb_46 = wdataMux_io_out_bits_wstrb_17;
  assign io_dram_wdata_bits_wstrb_47 = wdataMux_io_out_bits_wstrb_16;
  assign io_dram_wdata_bits_wstrb_48 = wdataMux_io_out_bits_wstrb_15;
  assign io_dram_wdata_bits_wstrb_49 = wdataMux_io_out_bits_wstrb_14;
  assign io_dram_wdata_bits_wstrb_50 = wdataMux_io_out_bits_wstrb_13;
  assign io_dram_wdata_bits_wstrb_51 = wdataMux_io_out_bits_wstrb_12;
  assign io_dram_wdata_bits_wstrb_52 = wdataMux_io_out_bits_wstrb_11;
  assign io_dram_wdata_bits_wstrb_53 = wdataMux_io_out_bits_wstrb_10;
  assign io_dram_wdata_bits_wstrb_54 = wdataMux_io_out_bits_wstrb_9;
  assign io_dram_wdata_bits_wstrb_55 = wdataMux_io_out_bits_wstrb_8;
  assign io_dram_wdata_bits_wstrb_56 = wdataMux_io_out_bits_wstrb_7;
  assign io_dram_wdata_bits_wstrb_57 = wdataMux_io_out_bits_wstrb_6;
  assign io_dram_wdata_bits_wstrb_58 = wdataMux_io_out_bits_wstrb_5;
  assign io_dram_wdata_bits_wstrb_59 = wdataMux_io_out_bits_wstrb_4;
  assign io_dram_wdata_bits_wstrb_60 = wdataMux_io_out_bits_wstrb_3;
  assign io_dram_wdata_bits_wstrb_61 = wdataMux_io_out_bits_wstrb_2;
  assign io_dram_wdata_bits_wstrb_62 = wdataMux_io_out_bits_wstrb_1;
  assign io_dram_wdata_bits_wstrb_63 = wdataMux_io_out_bits_wstrb_0;
  assign io_dram_rresp_ready = rrespReadyMux_io_out;
  assign io_dram_wresp_ready = wrespReadyMux_io_out;
  assign io_debugSignals_0 = FF_io_out[31:0];
  assign io_debugSignals_1 = {{26'd0}, FF_1_io_out};
  assign io_debugSignals_2 = FF_2_io_out[31:0];
  assign io_debugSignals_3 = FF_3_io_out;
  assign io_debugSignals_4 = {{31'd0}, FF_4_io_out};
  assign io_debugSignals_5 = {{16'd0}, FF_5_io_out};
  assign io_debugSignals_6 = Counter_io_out[31:0];
  assign io_debugSignals_7 = Counter_1_io_out[31:0];
  assign io_debugSignals_8 = Counter_2_io_out[31:0];
  assign io_debugSignals_9 = Counter_3_io_out[31:0];
  assign io_debugSignals_10 = Counter_4_io_out[31:0];
  assign io_debugSignals_11 = FF_6_io_out;
  assign io_debugSignals_12 = FF_7_io_out[31:0];
  assign io_debugSignals_13 = Counter_6_io_out[31:0];
  assign io_debugSignals_14 = Counter_7_io_out[31:0];
  assign io_debugSignals_15 = Counter_8_io_out[31:0];
  assign io_debugSignals_16 = cycleCount_io_out[31:0];
  assign io_debugSignals_17 = Counter_9_io_out[31:0];
  assign io_debugSignals_18 = Counter_10_io_out[31:0];
  assign io_debugSignals_19 = Counter_11_io_out[31:0];
  assign io_debugSignals_20 = Counter_13_io_out[31:0];
  assign io_debugSignals_21 = Counter_14_io_out[31:0];
  assign io_debugSignals_22 = Counter_12_io_out[31:0];
  assign io_debugSignals_23 = Counter_15_io_out[31:0];
  assign io_debugSignals_24 = Counter_17_io_out[31:0];
  assign io_debugSignals_25 = Counter_18_io_out[31:0];
  assign io_debugSignals_26 = Counter_16_io_out[31:0];
  assign io_debugSignals_27 = Counter_19_io_out[31:0];
  assign io_debugSignals_28 = Counter_20_io_out[31:0];
  assign io_debugSignals_29 = Counter_21_io_out[31:0];
  assign io_debugSignals_30 = Counter_22_io_out[31:0];
  assign io_debugSignals_31 = Counter_23_io_out[31:0];
  assign io_debugSignals_32 = Counter_24_io_out[31:0];
  assign io_debugSignals_33 = Counter_25_io_out[31:0];
  assign io_debugSignals_34 = Counter_26_io_out[31:0];
  assign io_debugSignals_35 = Counter_27_io_out[31:0];
  assign io_debugSignals_36 = Counter_28_io_out[31:0];
  assign io_debugSignals_37 = Counter_29_io_out[31:0];
  assign io_debugSignals_38 = Counter_30_io_out[31:0];
  assign io_debugSignals_39 = Counter_31_io_out[31:0];
  assign io_debugSignals_40 = Counter_32_io_out[31:0];
  assign io_debugSignals_41 = Counter_33_io_out[31:0];
  assign io_debugSignals_42 = Counter_34_io_out[31:0];
  assign io_debugSignals_43 = {{26'd0}, FF_9_io_out};
  assign io_debugSignals_44 = Counter_35_io_out[31:0];
  assign io_debugSignals_45 = Counter_36_io_out[31:0];
  assign io_debugSignals_46 = Counter_37_io_out[31:0];
  assign io_debugSignals_47 = Counter_38_io_out[31:0];
  assign io_debugSignals_48 = Counter_39_io_out[31:0];
  assign io_debugSignals_49 = Counter_40_io_out[31:0];
  assign io_debugSignals_50 = Counter_41_io_out[31:0];
  assign io_debugSignals_51 = Counter_42_io_out[31:0];
  assign io_debugSignals_52 = Counter_43_io_out[31:0];
  assign io_debugSignals_53 = Counter_44_io_out[31:0];
  assign io_debugSignals_54 = Counter_45_io_out[31:0];
  assign io_debugSignals_55 = Counter_46_io_out[31:0];
  assign io_debugSignals_56 = wdataCount_io_out[31:0];
  assign io_debugSignals_57 = Counter_47_io_out[31:0];
  assign io_debugSignals_58 = Counter_48_io_out[31:0];
  assign io_debugSignals_59 = Counter_49_io_out[31:0];
  assign io_debugSignals_60 = Counter_50_io_out[31:0];
  assign io_debugSignals_61 = Counter_51_io_out[31:0];
  assign io_debugSignals_62 = Counter_52_io_out[31:0];
  assign io_debugSignals_63 = Counter_53_io_out[31:0];
  assign io_debugSignals_64 = Counter_54_io_out[31:0];
  assign io_debugSignals_65 = Counter_55_io_out[31:0];
  assign io_debugSignals_66 = Counter_56_io_out[31:0];
  assign io_debugSignals_67 = Counter_57_io_out[31:0];
  assign io_debugSignals_68 = Counter_58_io_out[31:0];
  assign io_debugSignals_69 = Counter_59_io_out[31:0];
  assign io_debugSignals_70 = FF_10_io_out[31:0];
  assign io_debugSignals_71 = {{24'd0}, FF_11_io_out};
  assign io_debugSignals_72 = {{29'd0}, FF_12_io_out};
  assign io_debugSignals_73 = {{31'd0}, FF_13_io_out};
  assign io_debugSignals_74 = {{30'd0}, FF_14_io_out};
  assign io_debugSignals_75 = FF_15_io_out[31:0];
  assign io_debugSignals_76 = {{24'd0}, FF_16_io_out};
  assign io_debugSignals_77 = FF_17_io_out[31:0];
  assign io_debugSignals_78 = FF_18_io_out[31:0];
  assign io_debugSignals_79 = FF_19_io_out[31:0];
  assign io_debugSignals_80 = FF_20_io_out[31:0];
  assign io_debugSignals_81 = FF_21_io_out[31:0];
  assign io_debugSignals_82 = FF_22_io_out[31:0];
  assign io_debugSignals_83 = Counter_60_io_out[31:0];
  assign io_debugSignals_84 = Counter_61_io_out[31:0];
  assign io_debugSignals_85 = Counter_62_io_out[31:0];
  assign io_debugSignals_86 = Counter_63_io_out[31:0];
  assign io_debugSignals_87 = Counter_64_io_out[31:0];
  assign io_debugSignals_88 = Counter_65_io_out[31:0];
  assign io_debugSignals_89 = Counter_66_io_out[31:0];
  assign io_debugSignals_90 = Counter_67_io_out[31:0];
  assign io_debugSignals_91 = Counter_68_io_out[31:0];
  assign io_debugSignals_92 = Counter_69_io_out[31:0];
  assign io_debugSignals_93 = Counter_70_io_out[31:0];
  assign io_debugSignals_94 = Counter_71_io_out[31:0];
  assign io_debugSignals_95 = Counter_72_io_out[31:0];
  assign io_debugSignals_96 = FF_23_io_out[31:0];
  assign io_debugSignals_97 = {{24'd0}, FF_24_io_out};
  assign io_debugSignals_98 = {{29'd0}, FF_25_io_out};
  assign io_debugSignals_99 = {{30'd0}, FF_26_io_out};
  assign io_debugSignals_100 = FF_27_io_out[31:0];
  assign io_debugSignals_101 = {{24'd0}, FF_28_io_out};
  assign io_debugSignals_102 = FF_29_io_out[31:0];
  assign io_debugSignals_103 = FF_30_io_out[31:0];
  assign io_debugSignals_104 = FF_31_io_out[31:0];
  assign io_debugSignals_105 = FF_32_io_out[31:0];
  assign io_debugSignals_106 = FF_33_io_out[31:0];
  assign io_debugSignals_107 = FF_34_io_out[31:0];
  assign cmdArbiter_io_fifo_0_deq_0_addr = cmdFifos_0_io_deq_0_addr;
  assign cmdArbiter_io_fifo_0_deq_0_isWr = cmdFifos_0_io_deq_0_isWr;
  assign cmdArbiter_io_fifo_0_deq_0_size = cmdFifos_0_io_deq_0_size;
  assign cmdArbiter_io_fifo_0_full = cmdFifos_0_io_full;
  assign cmdArbiter_io_fifo_0_empty = cmdFifos_0_io_empty;
  assign cmdArbiter_io_fifo_0_almostEmpty = cmdFifos_0_io_almostEmpty;
  assign cmdArbiter_io_fifo_1_deq_0_addr = cmdFifos_1_io_deq_0_addr;
  assign cmdArbiter_io_fifo_1_deq_0_isWr = cmdFifos_1_io_deq_0_isWr;
  assign cmdArbiter_io_fifo_1_deq_0_size = cmdFifos_1_io_deq_0_size;
  assign cmdArbiter_io_fifo_1_empty = cmdFifos_1_io_empty;
  assign cmdArbiter_io_enq_0_0_addr = io_app_loads_0_cmd_bits_addr;
  assign cmdArbiter_io_enq_0_0_isWr = io_app_loads_0_cmd_bits_isWr;
  assign cmdArbiter_io_enq_0_0_size = io_app_loads_0_cmd_bits_size;
  assign cmdArbiter_io_enqVld_0 = io_app_loads_0_cmd_valid;
  assign cmdArbiter_io_deqVld = cmdDeqValidMux_io_out;
  assign cmdArbiter_clock = clock;
  assign cmdArbiter_reset = reset;
  assign cmdFifos_0_io_enq_0_addr = cmdArbiter_io_fifo_0_enq_0_addr;
  assign cmdFifos_0_io_enq_0_isWr = cmdArbiter_io_fifo_0_enq_0_isWr;
  assign cmdFifos_0_io_enq_0_size = cmdArbiter_io_fifo_0_enq_0_size;
  assign cmdFifos_0_io_enqVld = cmdArbiter_io_fifo_0_enqVld;
  assign cmdFifos_0_io_deqVld = cmdArbiter_io_fifo_0_deqVld;
  assign cmdFifos_0_clock = clock;
  assign cmdFifos_0_reset = reset;
  assign cmdFifos_1_io_enq_0_addr = 64'h0;
  assign cmdFifos_1_io_enq_0_isWr = 1'h0;
  assign cmdFifos_1_io_enq_0_size = 16'h0;
  assign cmdFifos_1_io_enqVld = 1'h0;
  assign cmdFifos_1_io_deqVld = cmdArbiter_io_fifo_1_deqVld;
  assign cmdFifos_1_clock = clock;
  assign cmdFifos_1_reset = reset;
  assign FF_io_in = _T_887;
  assign FF_io_init = 64'h175be;
  assign FF_io_reset = 1'h0;
  assign FF_io_enable = io_app_loads_0_cmd_valid;
  assign FF_clock = clock;
  assign FF_reset = reset;
  assign sizeCounter_io_max = _T_903;
  assign sizeCounter_io_stride = 16'h4000;
  assign sizeCounter_io_reset = 1'h0;
  assign sizeCounter_io_enable = _T_1197;
  assign sizeCounter_clock = clock;
  assign sizeCounter_reset = reset;
  assign cmdAddr_bits = _T_895;
  assign isSparseMux_io_ins_0 = 1'h0;
  assign isSparseMux_io_ins_1 = 1'h0;
  assign isSparseMux_io_sel = cmdArbiter_io_tag;
  assign burstCounter_io_max = _T_1231[15:0];
  assign burstCounter_io_stride = 16'h1;
  assign burstCounter_io_reset = io_reset;
  assign burstCounter_io_enable = _T_1235;
  assign burstCounter_clock = clock;
  assign burstCounter_reset = reset;
  assign burstTagCounter_io_reset = io_reset;
  assign burstTagCounter_io_enable = _T_1197;
  assign burstTagCounter_clock = clock;
  assign burstTagCounter_reset = reset;
  assign dramReadySeen = dramReadyFF_io_out;
  assign cmdCooldown_io_in = 1'h1;
  assign cmdCooldown_io_init = 1'h0;
  assign cmdCooldown_io_reset = _T_1249;
  assign cmdCooldown_io_enable = _T_1197;
  assign cmdCooldown_clock = clock;
  assign cmdCooldown_reset = reset;
  assign burstCounterDoneLatch_io_in = 1'h1;
  assign burstCounterDoneLatch_io_init = 1'h0;
  assign burstCounterDoneLatch_io_reset = _T_1229;
  assign burstCounterDoneLatch_io_enable = _T_1227;
  assign burstCounterDoneLatch_clock = clock;
  assign burstCounterDoneLatch_reset = reset;
  assign sizeCounterDoneLatch_io_in = 1'h1;
  assign sizeCounterDoneLatch_io_init = 1'h0;
  assign sizeCounterDoneLatch_io_reset = burstCounterDoneLatch_io_out;
  assign sizeCounterDoneLatch_io_enable = _T_908;
  assign sizeCounterDoneLatch_clock = clock;
  assign sizeCounterDoneLatch_reset = reset;
  assign rrespReadyMux_io_ins_0 = _T_1029;
  assign wdataMux_io_ins_0_valid = _T_1129;
  assign wdataMux_io_ins_0_bits_wdata_0 = denseStoreBuffers_0_io_deq_0;
  assign wdataMux_io_ins_0_bits_wdata_1 = denseStoreBuffers_0_io_deq_1;
  assign wdataMux_io_ins_0_bits_wdata_2 = denseStoreBuffers_0_io_deq_2;
  assign wdataMux_io_ins_0_bits_wdata_3 = denseStoreBuffers_0_io_deq_3;
  assign wdataMux_io_ins_0_bits_wdata_4 = denseStoreBuffers_0_io_deq_4;
  assign wdataMux_io_ins_0_bits_wdata_5 = denseStoreBuffers_0_io_deq_5;
  assign wdataMux_io_ins_0_bits_wdata_6 = denseStoreBuffers_0_io_deq_6;
  assign wdataMux_io_ins_0_bits_wdata_7 = denseStoreBuffers_0_io_deq_7;
  assign wdataMux_io_ins_0_bits_wdata_8 = denseStoreBuffers_0_io_deq_8;
  assign wdataMux_io_ins_0_bits_wdata_9 = denseStoreBuffers_0_io_deq_9;
  assign wdataMux_io_ins_0_bits_wdata_10 = denseStoreBuffers_0_io_deq_10;
  assign wdataMux_io_ins_0_bits_wdata_11 = denseStoreBuffers_0_io_deq_11;
  assign wdataMux_io_ins_0_bits_wdata_12 = denseStoreBuffers_0_io_deq_12;
  assign wdataMux_io_ins_0_bits_wdata_13 = denseStoreBuffers_0_io_deq_13;
  assign wdataMux_io_ins_0_bits_wdata_14 = denseStoreBuffers_0_io_deq_14;
  assign wdataMux_io_ins_0_bits_wdata_15 = denseStoreBuffers_0_io_deq_15;
  assign wdataMux_io_ins_0_bits_wstrb_0 = _T_1130;
  assign wdataMux_io_ins_0_bits_wstrb_1 = _T_1131;
  assign wdataMux_io_ins_0_bits_wstrb_2 = _T_1132;
  assign wdataMux_io_ins_0_bits_wstrb_3 = _T_1133;
  assign wdataMux_io_ins_0_bits_wstrb_4 = _T_1134;
  assign wdataMux_io_ins_0_bits_wstrb_5 = _T_1135;
  assign wdataMux_io_ins_0_bits_wstrb_6 = _T_1136;
  assign wdataMux_io_ins_0_bits_wstrb_7 = _T_1137;
  assign wdataMux_io_ins_0_bits_wstrb_8 = _T_1138;
  assign wdataMux_io_ins_0_bits_wstrb_9 = _T_1139;
  assign wdataMux_io_ins_0_bits_wstrb_10 = _T_1140;
  assign wdataMux_io_ins_0_bits_wstrb_11 = _T_1141;
  assign wdataMux_io_ins_0_bits_wstrb_12 = _T_1142;
  assign wdataMux_io_ins_0_bits_wstrb_13 = _T_1143;
  assign wdataMux_io_ins_0_bits_wstrb_14 = _T_1144;
  assign wdataMux_io_ins_0_bits_wstrb_15 = _T_1145;
  assign wdataMux_io_ins_0_bits_wstrb_16 = _T_1146;
  assign wdataMux_io_ins_0_bits_wstrb_17 = _T_1147;
  assign wdataMux_io_ins_0_bits_wstrb_18 = _T_1148;
  assign wdataMux_io_ins_0_bits_wstrb_19 = _T_1149;
  assign wdataMux_io_ins_0_bits_wstrb_20 = _T_1150;
  assign wdataMux_io_ins_0_bits_wstrb_21 = _T_1151;
  assign wdataMux_io_ins_0_bits_wstrb_22 = _T_1152;
  assign wdataMux_io_ins_0_bits_wstrb_23 = _T_1153;
  assign wdataMux_io_ins_0_bits_wstrb_24 = _T_1154;
  assign wdataMux_io_ins_0_bits_wstrb_25 = _T_1155;
  assign wdataMux_io_ins_0_bits_wstrb_26 = _T_1156;
  assign wdataMux_io_ins_0_bits_wstrb_27 = _T_1157;
  assign wdataMux_io_ins_0_bits_wstrb_28 = _T_1158;
  assign wdataMux_io_ins_0_bits_wstrb_29 = _T_1159;
  assign wdataMux_io_ins_0_bits_wstrb_30 = _T_1160;
  assign wdataMux_io_ins_0_bits_wstrb_31 = _T_1161;
  assign wdataMux_io_ins_0_bits_wstrb_32 = _T_1162;
  assign wdataMux_io_ins_0_bits_wstrb_33 = _T_1163;
  assign wdataMux_io_ins_0_bits_wstrb_34 = _T_1164;
  assign wdataMux_io_ins_0_bits_wstrb_35 = _T_1165;
  assign wdataMux_io_ins_0_bits_wstrb_36 = _T_1166;
  assign wdataMux_io_ins_0_bits_wstrb_37 = _T_1167;
  assign wdataMux_io_ins_0_bits_wstrb_38 = _T_1168;
  assign wdataMux_io_ins_0_bits_wstrb_39 = _T_1169;
  assign wdataMux_io_ins_0_bits_wstrb_40 = _T_1170;
  assign wdataMux_io_ins_0_bits_wstrb_41 = _T_1171;
  assign wdataMux_io_ins_0_bits_wstrb_42 = _T_1172;
  assign wdataMux_io_ins_0_bits_wstrb_43 = _T_1173;
  assign wdataMux_io_ins_0_bits_wstrb_44 = _T_1174;
  assign wdataMux_io_ins_0_bits_wstrb_45 = _T_1175;
  assign wdataMux_io_ins_0_bits_wstrb_46 = _T_1176;
  assign wdataMux_io_ins_0_bits_wstrb_47 = _T_1177;
  assign wdataMux_io_ins_0_bits_wstrb_48 = _T_1178;
  assign wdataMux_io_ins_0_bits_wstrb_49 = _T_1179;
  assign wdataMux_io_ins_0_bits_wstrb_50 = _T_1180;
  assign wdataMux_io_ins_0_bits_wstrb_51 = _T_1181;
  assign wdataMux_io_ins_0_bits_wstrb_52 = _T_1182;
  assign wdataMux_io_ins_0_bits_wstrb_53 = _T_1183;
  assign wdataMux_io_ins_0_bits_wstrb_54 = _T_1184;
  assign wdataMux_io_ins_0_bits_wstrb_55 = _T_1185;
  assign wdataMux_io_ins_0_bits_wstrb_56 = _T_1186;
  assign wdataMux_io_ins_0_bits_wstrb_57 = _T_1187;
  assign wdataMux_io_ins_0_bits_wstrb_58 = _T_1188;
  assign wdataMux_io_ins_0_bits_wstrb_59 = _T_1189;
  assign wdataMux_io_ins_0_bits_wstrb_60 = _T_1190;
  assign wdataMux_io_ins_0_bits_wstrb_61 = _T_1191;
  assign wdataMux_io_ins_0_bits_wstrb_62 = _T_1192;
  assign wdataMux_io_ins_0_bits_wstrb_63 = _T_1193;
  assign cmdDeqValidMux_io_ins_0 = sizeCounterDoneLatch_io_out;
  assign cmdDeqValidMux_io_ins_1 = _T_1109;
  assign cmdDeqValidMux_io_sel = cmdArbiter_io_tag;
  assign dramCmdMux_io_ins_0_valid = cmdRead;
  assign dramCmdMux_io_ins_0_bits_addr = _T_933;
  assign dramCmdMux_io_ins_0_bits_size = {{22'd0}, _T_949};
  assign dramCmdMux_io_ins_0_bits_isWr = cmdArbiter_io_deq_0_isWr;
  assign dramCmdMux_io_ins_0_bits_tag_uid = {{16'd0}, burstTagCounter_io_out};
  assign dramCmdMux_io_ins_0_bits_tag_streamId = _T_935_streamId;
  assign dramCmdMux_io_ins_1_valid = _T_1112;
  assign dramCmdMux_io_ins_1_bits_addr = _T_933;
  assign dramCmdMux_io_ins_1_bits_size = {{22'd0}, _T_983};
  assign dramCmdMux_io_ins_1_bits_isWr = cmdArbiter_io_deq_0_isWr;
  assign dramCmdMux_io_ins_1_bits_tag_uid = {{16'd0}, burstTagCounter_io_out};
  assign dramCmdMux_io_ins_1_bits_tag_streamId = _T_969_streamId;
  assign dramCmdMux_io_sel = cmdArbiter_io_tag;
  assign _T_935_streamId = {{5'd0}, cmdArbiter_io_tag};
  assign _T_937_bits = _T_943;
  assign FF_1_io_in = dramCmdMux_io_out_bits_tag_streamId;
  assign FF_1_io_enable = _T_951;
  assign FF_1_clock = clock;
  assign FF_1_reset = reset;
  assign FF_2_io_in = dramCmdMux_io_out_bits_addr;
  assign FF_2_io_init = 64'h2eb7e;
  assign FF_2_io_reset = 1'h0;
  assign FF_2_io_enable = _T_951;
  assign FF_2_clock = clock;
  assign FF_2_reset = reset;
  assign FF_3_io_in = dramCmdMux_io_out_bits_size;
  assign FF_3_io_enable = _T_951;
  assign FF_3_clock = clock;
  assign FF_3_reset = reset;
  assign _T_969_streamId = {{5'd0}, cmdArbiter_io_tag};
  assign _T_971_bits = _T_943;
  assign FF_4_io_in = cmdArbiter_io_tag;
  assign FF_4_io_init = 1'h0;
  assign FF_4_io_reset = 1'h0;
  assign FF_4_io_enable = cmdWrite;
  assign FF_4_clock = clock;
  assign FF_4_reset = reset;
  assign FF_5_io_in = cmdArbiter_io_deq_0_size;
  assign FF_5_io_enable = cmdWrite;
  assign FF_5_clock = clock;
  assign FF_5_reset = reset;
  assign wrespReadyMux_io_ins_0 = _T_1204;
  assign gatherLoadIssueMux_io_ins_0 = 1'h0;
  assign gatherLoadIssueMux_io_ins_1 = 1'h0;
  assign gatherLoadIssueMux_io_sel = cmdArbiter_io_tag;
  assign gatherLoadIssue_io_reset = io_reset;
  assign gatherLoadIssue_io_enable = gatherLoadIssueMux_io_out;
  assign gatherLoadIssue_clock = clock;
  assign gatherLoadIssue_reset = reset;
  assign gatherLoadSkipMux_io_ins_0 = 1'h0;
  assign gatherLoadSkipMux_io_ins_1 = 1'h0;
  assign gatherLoadSkipMux_io_sel = cmdArbiter_io_tag;
  assign gatherLoadSkip_io_reset = io_reset;
  assign gatherLoadSkip_io_enable = gatherLoadSkipMux_io_out;
  assign gatherLoadSkip_clock = clock;
  assign gatherLoadSkip_reset = reset;
  assign scatterLoadIssueMux_io_ins_0 = 1'h0;
  assign scatterLoadIssueMux_io_ins_1 = 1'h0;
  assign scatterLoadIssueMux_io_sel = cmdArbiter_io_tag;
  assign scatterLoadIssue_io_reset = io_reset;
  assign scatterLoadIssue_io_enable = scatterLoadIssueMux_io_out;
  assign scatterLoadIssue_clock = clock;
  assign scatterLoadIssue_reset = reset;
  assign scatterLoadSkipMux_io_ins_0 = 1'h0;
  assign scatterLoadSkipMux_io_ins_1 = 1'h0;
  assign scatterLoadSkipMux_io_sel = cmdArbiter_io_tag;
  assign scatterLoadSkip_io_reset = io_reset;
  assign scatterLoadSkip_io_enable = scatterLoadSkipMux_io_out;
  assign scatterLoadSkip_clock = clock;
  assign scatterLoadSkip_reset = reset;
  assign scatterStoreIssueMux_io_ins_0 = 1'h0;
  assign scatterStoreIssueMux_io_ins_1 = 1'h0;
  assign scatterStoreIssueMux_io_sel = cmdArbiter_io_tag;
  assign scatterStoreIssue_io_reset = io_reset;
  assign scatterStoreIssue_io_enable = scatterStoreIssueMux_io_out;
  assign scatterStoreIssue_clock = clock;
  assign scatterStoreIssue_reset = reset;
  assign scatterStoreSkipMux_io_ins_0 = 1'h0;
  assign scatterStoreSkipMux_io_ins_1 = 1'h0;
  assign scatterStoreSkipMux_io_sel = cmdArbiter_io_tag;
  assign scatterStoreSkip_io_reset = io_reset;
  assign scatterStoreSkip_io_enable = scatterStoreSkipMux_io_out;
  assign scatterStoreSkip_clock = clock;
  assign scatterStoreSkip_reset = reset;
  assign denseLoadBuffers_0_io_enq_0 = io_dram_rresp_bits_rdata_0;
  assign denseLoadBuffers_0_io_enq_1 = io_dram_rresp_bits_rdata_1;
  assign denseLoadBuffers_0_io_enq_2 = io_dram_rresp_bits_rdata_2;
  assign denseLoadBuffers_0_io_enq_3 = io_dram_rresp_bits_rdata_3;
  assign denseLoadBuffers_0_io_enq_4 = io_dram_rresp_bits_rdata_4;
  assign denseLoadBuffers_0_io_enq_5 = io_dram_rresp_bits_rdata_5;
  assign denseLoadBuffers_0_io_enq_6 = io_dram_rresp_bits_rdata_6;
  assign denseLoadBuffers_0_io_enq_7 = io_dram_rresp_bits_rdata_7;
  assign denseLoadBuffers_0_io_enq_8 = io_dram_rresp_bits_rdata_8;
  assign denseLoadBuffers_0_io_enq_9 = io_dram_rresp_bits_rdata_9;
  assign denseLoadBuffers_0_io_enq_10 = io_dram_rresp_bits_rdata_10;
  assign denseLoadBuffers_0_io_enq_11 = io_dram_rresp_bits_rdata_11;
  assign denseLoadBuffers_0_io_enq_12 = io_dram_rresp_bits_rdata_12;
  assign denseLoadBuffers_0_io_enq_13 = io_dram_rresp_bits_rdata_13;
  assign denseLoadBuffers_0_io_enq_14 = io_dram_rresp_bits_rdata_14;
  assign denseLoadBuffers_0_io_enq_15 = io_dram_rresp_bits_rdata_15;
  assign denseLoadBuffers_0_io_enqVld = _T_1028;
  assign denseLoadBuffers_0_io_deqVld = io_app_loads_0_rdata_ready;
  assign denseLoadBuffers_0_clock = clock;
  assign denseLoadBuffers_0_reset = reset;
  assign Counter_io_reset = io_reset;
  assign Counter_io_enable = denseLoadBuffers_0_io_enqVld;
  assign Counter_clock = clock;
  assign Counter_reset = reset;
  assign Counter_1_io_reset = io_reset;
  assign Counter_1_io_enable = _T_1031;
  assign Counter_1_clock = clock;
  assign Counter_1_reset = reset;
  assign Counter_2_io_reset = io_reset;
  assign Counter_2_io_enable = io_app_loads_0_rdata_ready;
  assign Counter_2_clock = clock;
  assign Counter_2_reset = reset;
  assign Counter_3_io_reset = io_reset;
  assign Counter_3_io_enable = _T_1046;
  assign Counter_3_clock = clock;
  assign Counter_3_reset = reset;
  assign Counter_4_io_reset = io_reset;
  assign Counter_4_io_enable = _T_1051;
  assign Counter_4_clock = clock;
  assign Counter_4_reset = reset;
  assign SRFF_io_input_set = denseLoadBuffers_0_io_deqVld;
  assign SRFF_io_input_reset = _T_1057;
  assign SRFF_io_input_asyn_reset = _T_1057;
  assign SRFF_clock = clock;
  assign SRFF_reset = reset;
  assign SRFF_1_io_input_set = denseLoadBuffers_0_io_enqVld;
  assign SRFF_1_io_input_reset = _T_1057;
  assign SRFF_1_io_input_asyn_reset = _T_1057;
  assign SRFF_1_clock = clock;
  assign SRFF_1_reset = reset;
  assign FF_6_io_in = denseLoadBuffers_0_io_deq_0;
  assign FF_6_io_enable = _T_1075;
  assign FF_6_clock = clock;
  assign FF_6_reset = reset;
  assign FF_7_io_in = _T_1105;
  assign FF_7_io_enable = _T_1090;
  assign FF_7_clock = clock;
  assign FF_7_reset = reset;
  assign denseStoreBuffers_0_io_enqVld = 1'h0;
  assign denseStoreBuffers_0_io_deqVld = _T_1123;
  assign denseStoreBuffers_0_clock = clock;
  assign denseStoreBuffers_0_reset = reset;
  assign Counter_5_io_max = FF_8_io_out;
  assign Counter_5_io_stride = 16'h4000;
  assign Counter_5_io_reset = 1'h0;
  assign Counter_5_io_enable = _T_1203;
  assign Counter_5_clock = clock;
  assign Counter_5_reset = reset;
  assign FF_8_io_in = cmdArbiter_io_deq_0_size;
  assign FF_8_io_enable = _T_1197;
  assign FF_8_clock = clock;
  assign FF_8_reset = reset;
  assign FIFOCounter_io_enqVld = Counter_5_io_done;
  assign FIFOCounter_clock = clock;
  assign FIFOCounter_reset = reset;
  assign Counter_6_io_reset = io_reset;
  assign Counter_6_io_enable = FIFOCounter_io_enqVld;
  assign Counter_6_clock = clock;
  assign Counter_6_reset = reset;
  assign Counter_7_io_reset = io_reset;
  assign Counter_7_io_enable = _T_1205;
  assign Counter_7_clock = clock;
  assign Counter_7_reset = reset;
  assign Counter_8_io_reset = io_reset;
  assign Counter_8_io_enable = 1'h0;
  assign Counter_8_clock = clock;
  assign Counter_8_reset = reset;
  assign burstCounterMaxLatch_io_in = io_dram_cmd_bits_size;
  assign burstCounterMaxLatch_io_enable = _T_1197;
  assign burstCounterMaxLatch_clock = clock;
  assign burstCounterMaxLatch_reset = reset;
  assign dramReadyFF_io_in = _T_1247;
  assign dramReadyFF_io_init = 1'h0;
  assign dramReadyFF_io_reset = 1'h0;
  assign dramReadyFF_io_enable = _T_1244;
  assign dramReadyFF_clock = clock;
  assign dramReadyFF_reset = reset;
  assign cycleCount_io_reset = io_reset;
  assign cycleCount_io_enable = io_enable;
  assign cycleCount_clock = clock;
  assign cycleCount_reset = reset;
  assign rdataEnqCount_io_reset = io_reset;
  assign rdataEnqCount_io_enable = _T_1261;
  assign rdataEnqCount_clock = clock;
  assign rdataEnqCount_reset = reset;
  assign wdataCount_io_reset = io_reset;
  assign wdataCount_io_enable = _T_1267;
  assign wdataCount_clock = clock;
  assign wdataCount_reset = reset;
  assign Counter_9_io_reset = io_reset;
  assign Counter_9_io_enable = _T_1273;
  assign Counter_9_clock = clock;
  assign Counter_9_reset = reset;
  assign Counter_10_io_reset = io_reset;
  assign Counter_10_io_enable = _T_1282;
  assign Counter_10_clock = clock;
  assign Counter_10_reset = reset;
  assign Counter_11_io_reset = io_reset;
  assign Counter_11_io_enable = _T_1290;
  assign Counter_11_clock = clock;
  assign Counter_11_reset = reset;
  assign Counter_12_io_reset = io_reset;
  assign Counter_12_io_enable = _T_1295;
  assign Counter_12_clock = clock;
  assign Counter_12_reset = reset;
  assign Counter_13_io_reset = io_reset;
  assign Counter_13_io_enable = _T_1301;
  assign Counter_13_clock = clock;
  assign Counter_13_reset = reset;
  assign Counter_14_io_reset = io_reset;
  assign Counter_14_io_enable = _T_1309;
  assign Counter_14_clock = clock;
  assign Counter_14_reset = reset;
  assign Counter_15_io_reset = io_reset;
  assign Counter_15_io_enable = _T_1316;
  assign Counter_15_clock = clock;
  assign Counter_15_reset = reset;
  assign Counter_16_io_reset = io_reset;
  assign Counter_16_io_enable = 1'h0;
  assign Counter_16_clock = clock;
  assign Counter_16_reset = reset;
  assign Counter_17_io_reset = io_reset;
  assign Counter_17_io_enable = 1'h0;
  assign Counter_17_clock = clock;
  assign Counter_17_reset = reset;
  assign Counter_18_io_reset = io_reset;
  assign Counter_18_io_enable = _T_1335;
  assign Counter_18_clock = clock;
  assign Counter_18_reset = reset;
  assign Counter_19_io_reset = io_reset;
  assign Counter_19_io_enable = _T_1261;
  assign Counter_19_clock = clock;
  assign Counter_19_reset = reset;
  assign Counter_20_io_reset = io_reset;
  assign Counter_20_io_enable = _T_1347;
  assign Counter_20_clock = clock;
  assign Counter_20_reset = reset;
  assign Counter_21_io_reset = io_reset;
  assign Counter_21_io_enable = _T_1354;
  assign Counter_21_clock = clock;
  assign Counter_21_reset = reset;
  assign Counter_22_io_reset = io_reset;
  assign Counter_22_io_enable = _T_1362;
  assign Counter_22_clock = clock;
  assign Counter_22_reset = reset;
  assign Counter_23_io_reset = io_reset;
  assign Counter_23_io_enable = _T_1367;
  assign Counter_23_clock = clock;
  assign Counter_23_reset = reset;
  assign Counter_24_io_reset = io_reset;
  assign Counter_24_io_enable = _T_1374;
  assign Counter_24_clock = clock;
  assign Counter_24_reset = reset;
  assign Counter_25_io_reset = io_reset;
  assign Counter_25_io_enable = _T_1381;
  assign Counter_25_clock = clock;
  assign Counter_25_reset = reset;
  assign Counter_26_io_reset = io_reset;
  assign Counter_26_io_enable = _T_1389;
  assign Counter_26_clock = clock;
  assign Counter_26_reset = reset;
  assign Counter_27_io_reset = io_reset;
  assign Counter_27_io_enable = denseLoadBuffers_0_io_full;
  assign Counter_27_clock = clock;
  assign Counter_27_reset = reset;
  assign Counter_28_io_reset = io_reset;
  assign Counter_28_io_enable = denseLoadBuffers_0_io_almostFull;
  assign Counter_28_clock = clock;
  assign Counter_28_reset = reset;
  assign Counter_29_io_reset = io_reset;
  assign Counter_29_io_enable = denseLoadBuffers_0_io_empty;
  assign Counter_29_clock = clock;
  assign Counter_29_reset = reset;
  assign Counter_30_io_reset = io_reset;
  assign Counter_30_io_enable = denseLoadBuffers_0_io_almostEmpty;
  assign Counter_30_clock = clock;
  assign Counter_30_reset = reset;
  assign Counter_31_io_reset = io_reset;
  assign Counter_31_io_enable = denseLoadBuffers_0_io_enqVld;
  assign Counter_31_clock = clock;
  assign Counter_31_reset = reset;
  assign Counter_32_io_reset = io_reset;
  assign Counter_32_io_enable = _T_1027;
  assign Counter_32_clock = clock;
  assign Counter_32_reset = reset;
  assign Counter_33_io_reset = io_reset;
  assign Counter_33_io_enable = io_dram_rresp_valid;
  assign Counter_33_clock = clock;
  assign Counter_33_reset = reset;
  assign Counter_34_io_reset = io_reset;
  assign Counter_34_io_enable = _T_1425;
  assign Counter_34_clock = clock;
  assign Counter_34_reset = reset;
  assign FF_9_io_in = io_dram_rresp_bits_tag_streamId;
  assign FF_9_io_enable = io_dram_rresp_valid;
  assign FF_9_clock = clock;
  assign FF_9_reset = reset;
  assign Counter_35_io_reset = io_reset;
  assign Counter_35_io_enable = denseStoreBuffers_0_io_enqVld;
  assign Counter_35_clock = clock;
  assign Counter_35_reset = reset;
  assign Counter_36_io_reset = io_reset;
  assign Counter_36_io_enable = _T_1194;
  assign Counter_36_clock = clock;
  assign Counter_36_reset = reset;
  assign Counter_37_io_reset = io_reset;
  assign Counter_37_io_enable = _T_1443;
  assign Counter_37_clock = clock;
  assign Counter_37_reset = reset;
  assign Counter_38_io_reset = io_reset;
  assign Counter_38_io_enable = _T_1448;
  assign Counter_38_clock = clock;
  assign Counter_38_reset = reset;
  assign Counter_39_io_reset = io_reset;
  assign Counter_39_io_enable = denseStoreBuffers_0_io_full;
  assign Counter_39_clock = clock;
  assign Counter_39_reset = reset;
  assign Counter_40_io_reset = io_reset;
  assign Counter_40_io_enable = denseStoreBuffers_0_io_almostFull;
  assign Counter_40_clock = clock;
  assign Counter_40_reset = reset;
  assign Counter_41_io_reset = io_reset;
  assign Counter_41_io_enable = denseStoreBuffers_0_io_empty;
  assign Counter_41_clock = clock;
  assign Counter_41_reset = reset;
  assign Counter_42_io_reset = io_reset;
  assign Counter_42_io_enable = denseStoreBuffers_0_io_almostEmpty;
  assign Counter_42_clock = clock;
  assign Counter_42_reset = reset;
  assign Counter_43_io_reset = io_reset;
  assign Counter_43_io_enable = _T_1469;
  assign Counter_43_clock = clock;
  assign Counter_43_reset = reset;
  assign Counter_44_io_reset = io_reset;
  assign Counter_44_io_enable = _T_1261;
  assign Counter_44_clock = clock;
  assign Counter_44_reset = reset;
  assign Counter_45_io_reset = io_reset;
  assign Counter_45_io_enable = _T_1480;
  assign Counter_45_clock = clock;
  assign Counter_45_reset = reset;
  assign Counter_46_io_reset = io_reset;
  assign Counter_46_io_enable = _T_1486;
  assign Counter_46_clock = clock;
  assign Counter_46_reset = reset;
  assign Counter_47_io_reset = io_reset;
  assign Counter_47_io_enable = io_TOP_AXI_ARVALID;
  assign Counter_47_clock = clock;
  assign Counter_47_reset = reset;
  assign Counter_48_io_reset = io_reset;
  assign Counter_48_io_enable = io_TOP_AXI_ARREADY;
  assign Counter_48_clock = clock;
  assign Counter_48_reset = reset;
  assign Counter_49_io_reset = io_reset;
  assign Counter_49_io_enable = _T_1499;
  assign Counter_49_clock = clock;
  assign Counter_49_reset = reset;
  assign Counter_50_io_reset = io_reset;
  assign Counter_50_io_enable = io_TOP_AXI_AWVALID;
  assign Counter_50_clock = clock;
  assign Counter_50_reset = reset;
  assign Counter_51_io_reset = io_reset;
  assign Counter_51_io_enable = _T_1508;
  assign Counter_51_clock = clock;
  assign Counter_51_reset = reset;
  assign Counter_52_io_reset = io_reset;
  assign Counter_52_io_enable = io_TOP_AXI_RVALID;
  assign Counter_52_clock = clock;
  assign Counter_52_reset = reset;
  assign Counter_53_io_reset = io_reset;
  assign Counter_53_io_enable = _T_1517;
  assign Counter_53_clock = clock;
  assign Counter_53_reset = reset;
  assign Counter_54_io_reset = io_reset;
  assign Counter_54_io_enable = io_TOP_AXI_WVALID;
  assign Counter_54_clock = clock;
  assign Counter_54_reset = reset;
  assign Counter_55_io_reset = io_reset;
  assign Counter_55_io_enable = _T_1526;
  assign Counter_55_clock = clock;
  assign Counter_55_reset = reset;
  assign Counter_56_io_reset = io_reset;
  assign Counter_56_io_enable = _T_1532;
  assign Counter_56_clock = clock;
  assign Counter_56_reset = reset;
  assign Counter_57_io_reset = io_reset;
  assign Counter_57_io_enable = _T_1531;
  assign Counter_57_clock = clock;
  assign Counter_57_reset = reset;
  assign Counter_58_io_reset = io_reset;
  assign Counter_58_io_enable = io_TOP_AXI_BVALID;
  assign Counter_58_clock = clock;
  assign Counter_58_reset = reset;
  assign Counter_59_io_reset = io_reset;
  assign Counter_59_io_enable = _T_1546;
  assign Counter_59_clock = clock;
  assign Counter_59_reset = reset;
  assign FF_10_io_in = io_TOP_AXI_ARADDR;
  assign FF_10_io_init = 64'h5d6fc6;
  assign FF_10_io_reset = 1'h0;
  assign FF_10_io_enable = _T_1551;
  assign FF_10_clock = clock;
  assign FF_10_reset = reset;
  assign FF_11_io_in = io_TOP_AXI_ARLEN;
  assign FF_11_io_enable = _T_1551;
  assign FF_11_clock = clock;
  assign FF_11_reset = reset;
  assign FF_12_io_in = io_TOP_AXI_ARSIZE;
  assign FF_12_io_enable = _T_1551;
  assign FF_12_clock = clock;
  assign FF_12_reset = reset;
  assign FF_13_io_in = io_TOP_AXI_ARID;
  assign FF_13_io_init = 1'h1;
  assign FF_13_io_reset = 1'h0;
  assign FF_13_io_enable = _T_1551;
  assign FF_13_clock = clock;
  assign FF_13_reset = reset;
  assign FF_14_io_in = io_TOP_AXI_ARBURST;
  assign FF_14_io_enable = _T_1551;
  assign FF_14_clock = clock;
  assign FF_14_reset = reset;
  assign FF_15_io_in = io_TOP_AXI_AWADDR;
  assign FF_15_io_init = 64'h5d6fcb;
  assign FF_15_io_reset = 1'h0;
  assign FF_15_io_enable = _T_1571;
  assign FF_15_clock = clock;
  assign FF_15_reset = reset;
  assign FF_16_io_in = io_TOP_AXI_AWLEN;
  assign FF_16_io_enable = _T_1571;
  assign FF_16_clock = clock;
  assign FF_16_reset = reset;
  assign FF_17_io_in = io_TOP_AXI_WDATA;
  assign FF_17_io_enable = _T_1579;
  assign FF_17_clock = clock;
  assign FF_17_reset = reset;
  assign FF_18_io_in = io_TOP_AXI_WSTRB;
  assign FF_18_io_init = 64'h5d6fce;
  assign FF_18_io_reset = 1'h0;
  assign FF_18_io_enable = _T_1579;
  assign FF_18_clock = clock;
  assign FF_18_reset = reset;
  assign FF_19_io_in = io_TOP_AXI_WDATA;
  assign FF_19_io_enable = _T_1590;
  assign FF_19_clock = clock;
  assign FF_19_reset = reset;
  assign FF_20_io_in = io_TOP_AXI_WSTRB;
  assign FF_20_io_init = 64'h5d6fd0;
  assign FF_20_io_reset = 1'h0;
  assign FF_20_io_enable = _T_1590;
  assign FF_20_clock = clock;
  assign FF_20_reset = reset;
  assign FF_21_io_in = io_TOP_AXI_WDATA;
  assign FF_21_io_enable = _T_1604;
  assign FF_21_clock = clock;
  assign FF_21_reset = reset;
  assign FF_22_io_in = io_TOP_AXI_WSTRB;
  assign FF_22_io_init = 64'h5d6fd2;
  assign FF_22_io_reset = 1'h0;
  assign FF_22_io_enable = _T_1604;
  assign FF_22_clock = clock;
  assign FF_22_reset = reset;
  assign Counter_60_io_reset = io_reset;
  assign Counter_60_io_enable = io_DWIDTH_AXI_ARVALID;
  assign Counter_60_clock = clock;
  assign Counter_60_reset = reset;
  assign Counter_61_io_reset = io_reset;
  assign Counter_61_io_enable = io_DWIDTH_AXI_ARREADY;
  assign Counter_61_clock = clock;
  assign Counter_61_reset = reset;
  assign Counter_62_io_reset = io_reset;
  assign Counter_62_io_enable = _T_1623;
  assign Counter_62_clock = clock;
  assign Counter_62_reset = reset;
  assign Counter_63_io_reset = io_reset;
  assign Counter_63_io_enable = io_DWIDTH_AXI_AWVALID;
  assign Counter_63_clock = clock;
  assign Counter_63_reset = reset;
  assign Counter_64_io_reset = io_reset;
  assign Counter_64_io_enable = _T_1632;
  assign Counter_64_clock = clock;
  assign Counter_64_reset = reset;
  assign Counter_65_io_reset = io_reset;
  assign Counter_65_io_enable = io_DWIDTH_AXI_RVALID;
  assign Counter_65_clock = clock;
  assign Counter_65_reset = reset;
  assign Counter_66_io_reset = io_reset;
  assign Counter_66_io_enable = _T_1641;
  assign Counter_66_clock = clock;
  assign Counter_66_reset = reset;
  assign Counter_67_io_reset = io_reset;
  assign Counter_67_io_enable = io_DWIDTH_AXI_WVALID;
  assign Counter_67_clock = clock;
  assign Counter_67_reset = reset;
  assign Counter_68_io_reset = io_reset;
  assign Counter_68_io_enable = _T_1650;
  assign Counter_68_clock = clock;
  assign Counter_68_reset = reset;
  assign Counter_69_io_reset = io_reset;
  assign Counter_69_io_enable = _T_1656;
  assign Counter_69_clock = clock;
  assign Counter_69_reset = reset;
  assign Counter_70_io_reset = io_reset;
  assign Counter_70_io_enable = _T_1655;
  assign Counter_70_clock = clock;
  assign Counter_70_reset = reset;
  assign Counter_71_io_reset = io_reset;
  assign Counter_71_io_enable = io_DWIDTH_AXI_BVALID;
  assign Counter_71_clock = clock;
  assign Counter_71_reset = reset;
  assign Counter_72_io_reset = io_reset;
  assign Counter_72_io_enable = _T_1670;
  assign Counter_72_clock = clock;
  assign Counter_72_reset = reset;
  assign FF_23_io_in = io_DWIDTH_AXI_ARADDR;
  assign FF_23_io_init = 64'h5d6fe0;
  assign FF_23_io_reset = 1'h0;
  assign FF_23_io_enable = _T_1675;
  assign FF_23_clock = clock;
  assign FF_23_reset = reset;
  assign FF_24_io_in = io_DWIDTH_AXI_ARLEN;
  assign FF_24_io_enable = _T_1675;
  assign FF_24_clock = clock;
  assign FF_24_reset = reset;
  assign FF_25_io_in = io_DWIDTH_AXI_ARSIZE;
  assign FF_25_io_enable = _T_1675;
  assign FF_25_clock = clock;
  assign FF_25_reset = reset;
  assign FF_26_io_in = io_DWIDTH_AXI_ARBURST;
  assign FF_26_io_enable = _T_1675;
  assign FF_26_clock = clock;
  assign FF_26_reset = reset;
  assign FF_27_io_in = io_DWIDTH_AXI_AWADDR;
  assign FF_27_io_init = 64'h5d6fe4;
  assign FF_27_io_reset = 1'h0;
  assign FF_27_io_enable = _T_1691;
  assign FF_27_clock = clock;
  assign FF_27_reset = reset;
  assign FF_28_io_in = io_DWIDTH_AXI_AWLEN;
  assign FF_28_io_enable = _T_1691;
  assign FF_28_clock = clock;
  assign FF_28_reset = reset;
  assign FF_29_io_in = io_DWIDTH_AXI_WDATA;
  assign FF_29_io_enable = _T_1699;
  assign FF_29_clock = clock;
  assign FF_29_reset = reset;
  assign FF_30_io_in = io_DWIDTH_AXI_WSTRB;
  assign FF_30_io_init = 64'h5d6fe7;
  assign FF_30_io_reset = 1'h0;
  assign FF_30_io_enable = _T_1699;
  assign FF_30_clock = clock;
  assign FF_30_reset = reset;
  assign FF_31_io_in = io_DWIDTH_AXI_WDATA;
  assign FF_31_io_enable = _T_1710;
  assign FF_31_clock = clock;
  assign FF_31_reset = reset;
  assign FF_32_io_in = io_DWIDTH_AXI_WSTRB;
  assign FF_32_io_init = 64'h5d6fe9;
  assign FF_32_io_reset = 1'h0;
  assign FF_32_io_enable = _T_1710;
  assign FF_32_clock = clock;
  assign FF_32_reset = reset;
  assign FF_33_io_in = io_DWIDTH_AXI_WDATA;
  assign FF_33_io_enable = _T_1724;
  assign FF_33_clock = clock;
  assign FF_33_reset = reset;
  assign FF_34_io_in = io_DWIDTH_AXI_WSTRB;
  assign FF_34_io_init = 64'h5d6feb;
  assign FF_34_io_reset = 1'h0;
  assign FF_34_io_enable = _T_1724;
  assign FF_34_clock = clock;
  assign FF_34_reset = reset;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_1068 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_1083 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_1068 <= 1'h0;
    end else begin
      _T_1068 <= _T_1065;
    end
    if (reset) begin
      _T_1083 <= 1'h0;
    end else begin
      _T_1083 <= _T_1080;
    end
  end
endmodule
module MAGCore_1(
  input         clock,
  input         reset,
  input         io_enable,
  input         io_reset,
  output        io_app_loads_0_cmd_ready,
  input         io_app_loads_0_cmd_valid,
  input  [63:0] io_app_loads_0_cmd_bits_addr,
  input         io_app_loads_0_cmd_bits_isWr,
  input  [15:0] io_app_loads_0_cmd_bits_size,
  input         io_app_loads_0_rdata_ready,
  output        io_app_loads_0_rdata_valid,
  output [31:0] io_app_loads_0_rdata_bits_0,
  input         io_dram_cmd_ready,
  output        io_dram_cmd_valid,
  output [63:0] io_dram_cmd_bits_addr,
  output [31:0] io_dram_cmd_bits_size,
  output        io_dram_cmd_bits_isWr,
  output [25:0] io_dram_cmd_bits_tag_uid,
  output [5:0]  io_dram_cmd_bits_tag_streamId,
  input         io_dram_wdata_ready,
  output        io_dram_wdata_valid,
  output [31:0] io_dram_wdata_bits_wdata_0,
  output [31:0] io_dram_wdata_bits_wdata_1,
  output [31:0] io_dram_wdata_bits_wdata_2,
  output [31:0] io_dram_wdata_bits_wdata_3,
  output [31:0] io_dram_wdata_bits_wdata_4,
  output [31:0] io_dram_wdata_bits_wdata_5,
  output [31:0] io_dram_wdata_bits_wdata_6,
  output [31:0] io_dram_wdata_bits_wdata_7,
  output [31:0] io_dram_wdata_bits_wdata_8,
  output [31:0] io_dram_wdata_bits_wdata_9,
  output [31:0] io_dram_wdata_bits_wdata_10,
  output [31:0] io_dram_wdata_bits_wdata_11,
  output [31:0] io_dram_wdata_bits_wdata_12,
  output [31:0] io_dram_wdata_bits_wdata_13,
  output [31:0] io_dram_wdata_bits_wdata_14,
  output [31:0] io_dram_wdata_bits_wdata_15,
  output        io_dram_wdata_bits_wstrb_0,
  output        io_dram_wdata_bits_wstrb_1,
  output        io_dram_wdata_bits_wstrb_2,
  output        io_dram_wdata_bits_wstrb_3,
  output        io_dram_wdata_bits_wstrb_4,
  output        io_dram_wdata_bits_wstrb_5,
  output        io_dram_wdata_bits_wstrb_6,
  output        io_dram_wdata_bits_wstrb_7,
  output        io_dram_wdata_bits_wstrb_8,
  output        io_dram_wdata_bits_wstrb_9,
  output        io_dram_wdata_bits_wstrb_10,
  output        io_dram_wdata_bits_wstrb_11,
  output        io_dram_wdata_bits_wstrb_12,
  output        io_dram_wdata_bits_wstrb_13,
  output        io_dram_wdata_bits_wstrb_14,
  output        io_dram_wdata_bits_wstrb_15,
  output        io_dram_wdata_bits_wstrb_16,
  output        io_dram_wdata_bits_wstrb_17,
  output        io_dram_wdata_bits_wstrb_18,
  output        io_dram_wdata_bits_wstrb_19,
  output        io_dram_wdata_bits_wstrb_20,
  output        io_dram_wdata_bits_wstrb_21,
  output        io_dram_wdata_bits_wstrb_22,
  output        io_dram_wdata_bits_wstrb_23,
  output        io_dram_wdata_bits_wstrb_24,
  output        io_dram_wdata_bits_wstrb_25,
  output        io_dram_wdata_bits_wstrb_26,
  output        io_dram_wdata_bits_wstrb_27,
  output        io_dram_wdata_bits_wstrb_28,
  output        io_dram_wdata_bits_wstrb_29,
  output        io_dram_wdata_bits_wstrb_30,
  output        io_dram_wdata_bits_wstrb_31,
  output        io_dram_wdata_bits_wstrb_32,
  output        io_dram_wdata_bits_wstrb_33,
  output        io_dram_wdata_bits_wstrb_34,
  output        io_dram_wdata_bits_wstrb_35,
  output        io_dram_wdata_bits_wstrb_36,
  output        io_dram_wdata_bits_wstrb_37,
  output        io_dram_wdata_bits_wstrb_38,
  output        io_dram_wdata_bits_wstrb_39,
  output        io_dram_wdata_bits_wstrb_40,
  output        io_dram_wdata_bits_wstrb_41,
  output        io_dram_wdata_bits_wstrb_42,
  output        io_dram_wdata_bits_wstrb_43,
  output        io_dram_wdata_bits_wstrb_44,
  output        io_dram_wdata_bits_wstrb_45,
  output        io_dram_wdata_bits_wstrb_46,
  output        io_dram_wdata_bits_wstrb_47,
  output        io_dram_wdata_bits_wstrb_48,
  output        io_dram_wdata_bits_wstrb_49,
  output        io_dram_wdata_bits_wstrb_50,
  output        io_dram_wdata_bits_wstrb_51,
  output        io_dram_wdata_bits_wstrb_52,
  output        io_dram_wdata_bits_wstrb_53,
  output        io_dram_wdata_bits_wstrb_54,
  output        io_dram_wdata_bits_wstrb_55,
  output        io_dram_wdata_bits_wstrb_56,
  output        io_dram_wdata_bits_wstrb_57,
  output        io_dram_wdata_bits_wstrb_58,
  output        io_dram_wdata_bits_wstrb_59,
  output        io_dram_wdata_bits_wstrb_60,
  output        io_dram_wdata_bits_wstrb_61,
  output        io_dram_wdata_bits_wstrb_62,
  output        io_dram_wdata_bits_wstrb_63,
  output        io_dram_rresp_ready,
  input         io_dram_rresp_valid,
  input  [31:0] io_dram_rresp_bits_rdata_0,
  input  [31:0] io_dram_rresp_bits_rdata_1,
  input  [31:0] io_dram_rresp_bits_rdata_2,
  input  [31:0] io_dram_rresp_bits_rdata_3,
  input  [31:0] io_dram_rresp_bits_rdata_4,
  input  [31:0] io_dram_rresp_bits_rdata_5,
  input  [31:0] io_dram_rresp_bits_rdata_6,
  input  [31:0] io_dram_rresp_bits_rdata_7,
  input  [31:0] io_dram_rresp_bits_rdata_8,
  input  [31:0] io_dram_rresp_bits_rdata_9,
  input  [31:0] io_dram_rresp_bits_rdata_10,
  input  [31:0] io_dram_rresp_bits_rdata_11,
  input  [31:0] io_dram_rresp_bits_rdata_12,
  input  [31:0] io_dram_rresp_bits_rdata_13,
  input  [31:0] io_dram_rresp_bits_rdata_14,
  input  [31:0] io_dram_rresp_bits_rdata_15,
  input  [5:0]  io_dram_rresp_bits_tag_streamId,
  output        io_dram_wresp_ready,
  input         io_dram_wresp_valid,
  input  [5:0]  io_dram_wresp_bits_tag_streamId
);
  wire  cmdArbiter_clock;
  wire  cmdArbiter_reset;
  wire [63:0] cmdArbiter_io_fifo_0_enq_0_addr;
  wire  cmdArbiter_io_fifo_0_enq_0_isWr;
  wire [15:0] cmdArbiter_io_fifo_0_enq_0_size;
  wire  cmdArbiter_io_fifo_0_enqVld;
  wire [63:0] cmdArbiter_io_fifo_0_deq_0_addr;
  wire  cmdArbiter_io_fifo_0_deq_0_isWr;
  wire [15:0] cmdArbiter_io_fifo_0_deq_0_size;
  wire  cmdArbiter_io_fifo_0_deqVld;
  wire  cmdArbiter_io_fifo_0_full;
  wire  cmdArbiter_io_fifo_0_empty;
  wire  cmdArbiter_io_fifo_0_almostEmpty;
  wire [63:0] cmdArbiter_io_fifo_1_deq_0_addr;
  wire  cmdArbiter_io_fifo_1_deq_0_isWr;
  wire [15:0] cmdArbiter_io_fifo_1_deq_0_size;
  wire  cmdArbiter_io_fifo_1_deqVld;
  wire  cmdArbiter_io_fifo_1_empty;
  wire [63:0] cmdArbiter_io_enq_0_0_addr;
  wire  cmdArbiter_io_enq_0_0_isWr;
  wire [15:0] cmdArbiter_io_enq_0_0_size;
  wire  cmdArbiter_io_enqVld_0;
  wire  cmdArbiter_io_full_0;
  wire [63:0] cmdArbiter_io_deq_0_addr;
  wire  cmdArbiter_io_deq_0_isWr;
  wire [15:0] cmdArbiter_io_deq_0_size;
  wire  cmdArbiter_io_deqVld;
  wire  cmdArbiter_io_deqReady;
  wire  cmdArbiter_io_empty;
  wire  cmdArbiter_io_tag;
  wire  cmdFifos_0_clock;
  wire  cmdFifos_0_reset;
  wire [63:0] cmdFifos_0_io_enq_0_addr;
  wire  cmdFifos_0_io_enq_0_isWr;
  wire [15:0] cmdFifos_0_io_enq_0_size;
  wire  cmdFifos_0_io_enqVld;
  wire [63:0] cmdFifos_0_io_deq_0_addr;
  wire  cmdFifos_0_io_deq_0_isWr;
  wire [15:0] cmdFifos_0_io_deq_0_size;
  wire  cmdFifos_0_io_deqVld;
  wire  cmdFifos_0_io_full;
  wire  cmdFifos_0_io_empty;
  wire  cmdFifos_0_io_almostEmpty;
  wire  cmdFifos_1_clock;
  wire  cmdFifos_1_reset;
  wire [63:0] cmdFifos_1_io_enq_0_addr;
  wire  cmdFifos_1_io_enq_0_isWr;
  wire [15:0] cmdFifos_1_io_enq_0_size;
  wire  cmdFifos_1_io_enqVld;
  wire [63:0] cmdFifos_1_io_deq_0_addr;
  wire  cmdFifos_1_io_deq_0_isWr;
  wire [15:0] cmdFifos_1_io_deq_0_size;
  wire  cmdFifos_1_io_deqVld;
  wire  cmdFifos_1_io_full;
  wire  cmdFifos_1_io_empty;
  wire  cmdFifos_1_io_almostEmpty;
  wire [31:0] _T_886;
  wire [63:0] _T_887;
  wire  FF_clock;
  wire  FF_reset;
  wire [63:0] FF_io_in;
  wire [63:0] FF_io_init;
  wire  FF_io_reset;
  wire [63:0] FF_io_out;
  wire  FF_io_enable;
  wire  sizeCounter_clock;
  wire  sizeCounter_reset;
  wire [15:0] sizeCounter_io_max;
  wire [15:0] sizeCounter_io_stride;
  wire [15:0] sizeCounter_io_out;
  wire  sizeCounter_io_last;
  wire  sizeCounter_io_reset;
  wire  sizeCounter_io_enable;
  wire  sizeCounter_io_done;
  wire  _T_891;
  wire [63:0] cmdAddr_bits;
  wire [63:0] _GEN_0;
  wire [64:0] _T_894;
  wire [63:0] _T_895;
  wire  _T_896;
  wire  _T_897;
  wire  cmdRead;
  wire  cmdWrite;
  wire  isSparseMux_io_ins_0;
  wire  isSparseMux_io_ins_1;
  wire  isSparseMux_io_sel;
  wire  isSparseMux_io_out;
  wire  burstCounter_clock;
  wire  burstCounter_reset;
  wire [15:0] burstCounter_io_max;
  wire [15:0] burstCounter_io_stride;
  wire [15:0] burstCounter_io_out;
  wire  burstCounter_io_last;
  wire  burstCounter_io_reset;
  wire  burstCounter_io_enable;
  wire  burstCounter_io_done;
  wire  burstTagCounter_clock;
  wire  burstTagCounter_reset;
  wire [9:0] burstTagCounter_io_out;
  wire  burstTagCounter_io_reset;
  wire  burstTagCounter_io_enable;
  wire  dramReadySeen;
  wire [15:0] _T_903;
  wire  cmdCooldown_clock;
  wire  cmdCooldown_reset;
  wire  cmdCooldown_io_in;
  wire  cmdCooldown_io_init;
  wire  cmdCooldown_io_reset;
  wire  cmdCooldown_io_out;
  wire  cmdCooldown_io_enable;
  wire  burstCounterDoneLatch_clock;
  wire  burstCounterDoneLatch_reset;
  wire  burstCounterDoneLatch_io_in;
  wire  burstCounterDoneLatch_io_init;
  wire  burstCounterDoneLatch_io_reset;
  wire  burstCounterDoneLatch_io_out;
  wire  burstCounterDoneLatch_io_enable;
  wire  sizeCounterDoneLatch_clock;
  wire  sizeCounterDoneLatch_reset;
  wire  sizeCounterDoneLatch_io_in;
  wire  sizeCounterDoneLatch_io_init;
  wire  sizeCounterDoneLatch_io_reset;
  wire  sizeCounterDoneLatch_io_out;
  wire  sizeCounterDoneLatch_io_enable;
  wire  _T_908;
  wire  rrespReadyMux_io_ins_0;
  wire  rrespReadyMux_io_out;
  wire  wdataMux_io_ins_0_valid;
  wire [31:0] wdataMux_io_ins_0_bits_wdata_0;
  wire [31:0] wdataMux_io_ins_0_bits_wdata_1;
  wire [31:0] wdataMux_io_ins_0_bits_wdata_2;
  wire [31:0] wdataMux_io_ins_0_bits_wdata_3;
  wire [31:0] wdataMux_io_ins_0_bits_wdata_4;
  wire [31:0] wdataMux_io_ins_0_bits_wdata_5;
  wire [31:0] wdataMux_io_ins_0_bits_wdata_6;
  wire [31:0] wdataMux_io_ins_0_bits_wdata_7;
  wire [31:0] wdataMux_io_ins_0_bits_wdata_8;
  wire [31:0] wdataMux_io_ins_0_bits_wdata_9;
  wire [31:0] wdataMux_io_ins_0_bits_wdata_10;
  wire [31:0] wdataMux_io_ins_0_bits_wdata_11;
  wire [31:0] wdataMux_io_ins_0_bits_wdata_12;
  wire [31:0] wdataMux_io_ins_0_bits_wdata_13;
  wire [31:0] wdataMux_io_ins_0_bits_wdata_14;
  wire [31:0] wdataMux_io_ins_0_bits_wdata_15;
  wire  wdataMux_io_ins_0_bits_wstrb_0;
  wire  wdataMux_io_ins_0_bits_wstrb_1;
  wire  wdataMux_io_ins_0_bits_wstrb_2;
  wire  wdataMux_io_ins_0_bits_wstrb_3;
  wire  wdataMux_io_ins_0_bits_wstrb_4;
  wire  wdataMux_io_ins_0_bits_wstrb_5;
  wire  wdataMux_io_ins_0_bits_wstrb_6;
  wire  wdataMux_io_ins_0_bits_wstrb_7;
  wire  wdataMux_io_ins_0_bits_wstrb_8;
  wire  wdataMux_io_ins_0_bits_wstrb_9;
  wire  wdataMux_io_ins_0_bits_wstrb_10;
  wire  wdataMux_io_ins_0_bits_wstrb_11;
  wire  wdataMux_io_ins_0_bits_wstrb_12;
  wire  wdataMux_io_ins_0_bits_wstrb_13;
  wire  wdataMux_io_ins_0_bits_wstrb_14;
  wire  wdataMux_io_ins_0_bits_wstrb_15;
  wire  wdataMux_io_ins_0_bits_wstrb_16;
  wire  wdataMux_io_ins_0_bits_wstrb_17;
  wire  wdataMux_io_ins_0_bits_wstrb_18;
  wire  wdataMux_io_ins_0_bits_wstrb_19;
  wire  wdataMux_io_ins_0_bits_wstrb_20;
  wire  wdataMux_io_ins_0_bits_wstrb_21;
  wire  wdataMux_io_ins_0_bits_wstrb_22;
  wire  wdataMux_io_ins_0_bits_wstrb_23;
  wire  wdataMux_io_ins_0_bits_wstrb_24;
  wire  wdataMux_io_ins_0_bits_wstrb_25;
  wire  wdataMux_io_ins_0_bits_wstrb_26;
  wire  wdataMux_io_ins_0_bits_wstrb_27;
  wire  wdataMux_io_ins_0_bits_wstrb_28;
  wire  wdataMux_io_ins_0_bits_wstrb_29;
  wire  wdataMux_io_ins_0_bits_wstrb_30;
  wire  wdataMux_io_ins_0_bits_wstrb_31;
  wire  wdataMux_io_ins_0_bits_wstrb_32;
  wire  wdataMux_io_ins_0_bits_wstrb_33;
  wire  wdataMux_io_ins_0_bits_wstrb_34;
  wire  wdataMux_io_ins_0_bits_wstrb_35;
  wire  wdataMux_io_ins_0_bits_wstrb_36;
  wire  wdataMux_io_ins_0_bits_wstrb_37;
  wire  wdataMux_io_ins_0_bits_wstrb_38;
  wire  wdataMux_io_ins_0_bits_wstrb_39;
  wire  wdataMux_io_ins_0_bits_wstrb_40;
  wire  wdataMux_io_ins_0_bits_wstrb_41;
  wire  wdataMux_io_ins_0_bits_wstrb_42;
  wire  wdataMux_io_ins_0_bits_wstrb_43;
  wire  wdataMux_io_ins_0_bits_wstrb_44;
  wire  wdataMux_io_ins_0_bits_wstrb_45;
  wire  wdataMux_io_ins_0_bits_wstrb_46;
  wire  wdataMux_io_ins_0_bits_wstrb_47;
  wire  wdataMux_io_ins_0_bits_wstrb_48;
  wire  wdataMux_io_ins_0_bits_wstrb_49;
  wire  wdataMux_io_ins_0_bits_wstrb_50;
  wire  wdataMux_io_ins_0_bits_wstrb_51;
  wire  wdataMux_io_ins_0_bits_wstrb_52;
  wire  wdataMux_io_ins_0_bits_wstrb_53;
  wire  wdataMux_io_ins_0_bits_wstrb_54;
  wire  wdataMux_io_ins_0_bits_wstrb_55;
  wire  wdataMux_io_ins_0_bits_wstrb_56;
  wire  wdataMux_io_ins_0_bits_wstrb_57;
  wire  wdataMux_io_ins_0_bits_wstrb_58;
  wire  wdataMux_io_ins_0_bits_wstrb_59;
  wire  wdataMux_io_ins_0_bits_wstrb_60;
  wire  wdataMux_io_ins_0_bits_wstrb_61;
  wire  wdataMux_io_ins_0_bits_wstrb_62;
  wire  wdataMux_io_ins_0_bits_wstrb_63;
  wire  wdataMux_io_out_valid;
  wire [31:0] wdataMux_io_out_bits_wdata_0;
  wire [31:0] wdataMux_io_out_bits_wdata_1;
  wire [31:0] wdataMux_io_out_bits_wdata_2;
  wire [31:0] wdataMux_io_out_bits_wdata_3;
  wire [31:0] wdataMux_io_out_bits_wdata_4;
  wire [31:0] wdataMux_io_out_bits_wdata_5;
  wire [31:0] wdataMux_io_out_bits_wdata_6;
  wire [31:0] wdataMux_io_out_bits_wdata_7;
  wire [31:0] wdataMux_io_out_bits_wdata_8;
  wire [31:0] wdataMux_io_out_bits_wdata_9;
  wire [31:0] wdataMux_io_out_bits_wdata_10;
  wire [31:0] wdataMux_io_out_bits_wdata_11;
  wire [31:0] wdataMux_io_out_bits_wdata_12;
  wire [31:0] wdataMux_io_out_bits_wdata_13;
  wire [31:0] wdataMux_io_out_bits_wdata_14;
  wire [31:0] wdataMux_io_out_bits_wdata_15;
  wire  wdataMux_io_out_bits_wstrb_0;
  wire  wdataMux_io_out_bits_wstrb_1;
  wire  wdataMux_io_out_bits_wstrb_2;
  wire  wdataMux_io_out_bits_wstrb_3;
  wire  wdataMux_io_out_bits_wstrb_4;
  wire  wdataMux_io_out_bits_wstrb_5;
  wire  wdataMux_io_out_bits_wstrb_6;
  wire  wdataMux_io_out_bits_wstrb_7;
  wire  wdataMux_io_out_bits_wstrb_8;
  wire  wdataMux_io_out_bits_wstrb_9;
  wire  wdataMux_io_out_bits_wstrb_10;
  wire  wdataMux_io_out_bits_wstrb_11;
  wire  wdataMux_io_out_bits_wstrb_12;
  wire  wdataMux_io_out_bits_wstrb_13;
  wire  wdataMux_io_out_bits_wstrb_14;
  wire  wdataMux_io_out_bits_wstrb_15;
  wire  wdataMux_io_out_bits_wstrb_16;
  wire  wdataMux_io_out_bits_wstrb_17;
  wire  wdataMux_io_out_bits_wstrb_18;
  wire  wdataMux_io_out_bits_wstrb_19;
  wire  wdataMux_io_out_bits_wstrb_20;
  wire  wdataMux_io_out_bits_wstrb_21;
  wire  wdataMux_io_out_bits_wstrb_22;
  wire  wdataMux_io_out_bits_wstrb_23;
  wire  wdataMux_io_out_bits_wstrb_24;
  wire  wdataMux_io_out_bits_wstrb_25;
  wire  wdataMux_io_out_bits_wstrb_26;
  wire  wdataMux_io_out_bits_wstrb_27;
  wire  wdataMux_io_out_bits_wstrb_28;
  wire  wdataMux_io_out_bits_wstrb_29;
  wire  wdataMux_io_out_bits_wstrb_30;
  wire  wdataMux_io_out_bits_wstrb_31;
  wire  wdataMux_io_out_bits_wstrb_32;
  wire  wdataMux_io_out_bits_wstrb_33;
  wire  wdataMux_io_out_bits_wstrb_34;
  wire  wdataMux_io_out_bits_wstrb_35;
  wire  wdataMux_io_out_bits_wstrb_36;
  wire  wdataMux_io_out_bits_wstrb_37;
  wire  wdataMux_io_out_bits_wstrb_38;
  wire  wdataMux_io_out_bits_wstrb_39;
  wire  wdataMux_io_out_bits_wstrb_40;
  wire  wdataMux_io_out_bits_wstrb_41;
  wire  wdataMux_io_out_bits_wstrb_42;
  wire  wdataMux_io_out_bits_wstrb_43;
  wire  wdataMux_io_out_bits_wstrb_44;
  wire  wdataMux_io_out_bits_wstrb_45;
  wire  wdataMux_io_out_bits_wstrb_46;
  wire  wdataMux_io_out_bits_wstrb_47;
  wire  wdataMux_io_out_bits_wstrb_48;
  wire  wdataMux_io_out_bits_wstrb_49;
  wire  wdataMux_io_out_bits_wstrb_50;
  wire  wdataMux_io_out_bits_wstrb_51;
  wire  wdataMux_io_out_bits_wstrb_52;
  wire  wdataMux_io_out_bits_wstrb_53;
  wire  wdataMux_io_out_bits_wstrb_54;
  wire  wdataMux_io_out_bits_wstrb_55;
  wire  wdataMux_io_out_bits_wstrb_56;
  wire  wdataMux_io_out_bits_wstrb_57;
  wire  wdataMux_io_out_bits_wstrb_58;
  wire  wdataMux_io_out_bits_wstrb_59;
  wire  wdataMux_io_out_bits_wstrb_60;
  wire  wdataMux_io_out_bits_wstrb_61;
  wire  wdataMux_io_out_bits_wstrb_62;
  wire  wdataMux_io_out_bits_wstrb_63;
  wire  cmdDeqValidMux_io_ins_0;
  wire  cmdDeqValidMux_io_ins_1;
  wire  cmdDeqValidMux_io_sel;
  wire  cmdDeqValidMux_io_out;
  wire  dramCmdMux_io_ins_0_valid;
  wire [63:0] dramCmdMux_io_ins_0_bits_addr;
  wire [31:0] dramCmdMux_io_ins_0_bits_size;
  wire  dramCmdMux_io_ins_0_bits_isWr;
  wire [25:0] dramCmdMux_io_ins_0_bits_tag_uid;
  wire [5:0] dramCmdMux_io_ins_0_bits_tag_streamId;
  wire  dramCmdMux_io_ins_1_valid;
  wire [63:0] dramCmdMux_io_ins_1_bits_addr;
  wire [31:0] dramCmdMux_io_ins_1_bits_size;
  wire  dramCmdMux_io_ins_1_bits_isWr;
  wire [25:0] dramCmdMux_io_ins_1_bits_tag_uid;
  wire [5:0] dramCmdMux_io_ins_1_bits_tag_streamId;
  wire  dramCmdMux_io_sel;
  wire  dramCmdMux_io_out_valid;
  wire [63:0] dramCmdMux_io_out_bits_addr;
  wire [31:0] dramCmdMux_io_out_bits_size;
  wire  dramCmdMux_io_out_bits_isWr;
  wire [25:0] dramCmdMux_io_out_bits_tag_uid;
  wire [5:0] dramCmdMux_io_out_bits_tag_streamId;
  wire [57:0] _T_931;
  wire [63:0] _T_933;
  wire [5:0] _T_935_streamId;
  wire [15:0] _T_937_bits;
  wire [16:0] _T_938;
  wire [16:0] _T_939;
  wire [15:0] _T_940;
  wire [15:0] _T_942;
  wire [15:0] _T_943;
  wire [9:0] _T_944;
  wire [5:0] _T_945;
  wire  _T_947;
  wire [9:0] _GEN_2;
  wire [10:0] _T_948;
  wire [9:0] _T_949;
  wire  _T_950;
  wire  _T_951;
  wire  FF_1_clock;
  wire  FF_1_reset;
  wire [5:0] FF_1_io_in;
  wire [5:0] FF_1_io_out;
  wire  FF_1_io_enable;
  wire  FF_2_clock;
  wire  FF_2_reset;
  wire [63:0] FF_2_io_in;
  wire [63:0] FF_2_io_init;
  wire  FF_2_io_reset;
  wire [63:0] FF_2_io_out;
  wire  FF_2_io_enable;
  wire  FF_3_clock;
  wire  FF_3_reset;
  wire [31:0] FF_3_io_in;
  wire [31:0] FF_3_io_out;
  wire  FF_3_io_enable;
  wire [5:0] _T_969_streamId;
  wire [15:0] _T_971_bits;
  wire [9:0] _T_978;
  wire [5:0] _T_979;
  wire  _T_981;
  wire [9:0] _GEN_3;
  wire [10:0] _T_982;
  wire [9:0] _T_983;
  wire  FF_4_clock;
  wire  FF_4_reset;
  wire  FF_4_io_in;
  wire  FF_4_io_init;
  wire  FF_4_io_reset;
  wire  FF_4_io_out;
  wire  FF_4_io_enable;
  wire  FF_5_clock;
  wire  FF_5_reset;
  wire [15:0] FF_5_io_in;
  wire [15:0] FF_5_io_out;
  wire  FF_5_io_enable;
  wire  wrespReadyMux_io_ins_0;
  wire  wrespReadyMux_io_out;
  wire  gatherLoadIssueMux_io_ins_0;
  wire  gatherLoadIssueMux_io_ins_1;
  wire  gatherLoadIssueMux_io_sel;
  wire  gatherLoadIssueMux_io_out;
  wire  gatherLoadIssue_clock;
  wire  gatherLoadIssue_reset;
  wire [63:0] gatherLoadIssue_io_out;
  wire  gatherLoadIssue_io_reset;
  wire  gatherLoadIssue_io_enable;
  wire  gatherLoadSkipMux_io_ins_0;
  wire  gatherLoadSkipMux_io_ins_1;
  wire  gatherLoadSkipMux_io_sel;
  wire  gatherLoadSkipMux_io_out;
  wire  gatherLoadSkip_clock;
  wire  gatherLoadSkip_reset;
  wire [63:0] gatherLoadSkip_io_out;
  wire  gatherLoadSkip_io_reset;
  wire  gatherLoadSkip_io_enable;
  wire  scatterLoadIssueMux_io_ins_0;
  wire  scatterLoadIssueMux_io_ins_1;
  wire  scatterLoadIssueMux_io_sel;
  wire  scatterLoadIssueMux_io_out;
  wire  scatterLoadIssue_clock;
  wire  scatterLoadIssue_reset;
  wire [63:0] scatterLoadIssue_io_out;
  wire  scatterLoadIssue_io_reset;
  wire  scatterLoadIssue_io_enable;
  wire  scatterLoadSkipMux_io_ins_0;
  wire  scatterLoadSkipMux_io_ins_1;
  wire  scatterLoadSkipMux_io_sel;
  wire  scatterLoadSkipMux_io_out;
  wire  scatterLoadSkip_clock;
  wire  scatterLoadSkip_reset;
  wire [63:0] scatterLoadSkip_io_out;
  wire  scatterLoadSkip_io_reset;
  wire  scatterLoadSkip_io_enable;
  wire  scatterStoreIssueMux_io_ins_0;
  wire  scatterStoreIssueMux_io_ins_1;
  wire  scatterStoreIssueMux_io_sel;
  wire  scatterStoreIssueMux_io_out;
  wire  scatterStoreIssue_clock;
  wire  scatterStoreIssue_reset;
  wire [63:0] scatterStoreIssue_io_out;
  wire  scatterStoreIssue_io_reset;
  wire  scatterStoreIssue_io_enable;
  wire  scatterStoreSkipMux_io_ins_0;
  wire  scatterStoreSkipMux_io_ins_1;
  wire  scatterStoreSkipMux_io_sel;
  wire  scatterStoreSkipMux_io_out;
  wire  scatterStoreSkip_clock;
  wire  scatterStoreSkip_reset;
  wire [63:0] scatterStoreSkip_io_out;
  wire  scatterStoreSkip_io_reset;
  wire  scatterStoreSkip_io_enable;
  wire  denseLoadBuffers_0_clock;
  wire  denseLoadBuffers_0_reset;
  wire [31:0] denseLoadBuffers_0_io_enq_0;
  wire [31:0] denseLoadBuffers_0_io_enq_1;
  wire [31:0] denseLoadBuffers_0_io_enq_2;
  wire [31:0] denseLoadBuffers_0_io_enq_3;
  wire [31:0] denseLoadBuffers_0_io_enq_4;
  wire [31:0] denseLoadBuffers_0_io_enq_5;
  wire [31:0] denseLoadBuffers_0_io_enq_6;
  wire [31:0] denseLoadBuffers_0_io_enq_7;
  wire [31:0] denseLoadBuffers_0_io_enq_8;
  wire [31:0] denseLoadBuffers_0_io_enq_9;
  wire [31:0] denseLoadBuffers_0_io_enq_10;
  wire [31:0] denseLoadBuffers_0_io_enq_11;
  wire [31:0] denseLoadBuffers_0_io_enq_12;
  wire [31:0] denseLoadBuffers_0_io_enq_13;
  wire [31:0] denseLoadBuffers_0_io_enq_14;
  wire [31:0] denseLoadBuffers_0_io_enq_15;
  wire  denseLoadBuffers_0_io_enqVld;
  wire [31:0] denseLoadBuffers_0_io_deq_0;
  wire  denseLoadBuffers_0_io_deqVld;
  wire  denseLoadBuffers_0_io_full;
  wire  denseLoadBuffers_0_io_empty;
  wire  denseLoadBuffers_0_io_almostEmpty;
  wire  denseLoadBuffers_0_io_almostFull;
  wire  _T_1027;
  wire  _T_1028;
  wire  _T_1029;
  wire  _T_1031;
  wire  Counter_clock;
  wire  Counter_reset;
  wire [63:0] Counter_io_out;
  wire  Counter_io_reset;
  wire  Counter_io_enable;
  wire  Counter_1_clock;
  wire  Counter_1_reset;
  wire [63:0] Counter_1_io_out;
  wire  Counter_1_io_reset;
  wire  Counter_1_io_enable;
  wire  Counter_2_clock;
  wire  Counter_2_reset;
  wire [63:0] Counter_2_io_out;
  wire  Counter_2_io_reset;
  wire  Counter_2_io_enable;
  wire  _T_1046;
  wire  Counter_3_clock;
  wire  Counter_3_reset;
  wire [63:0] Counter_3_io_out;
  wire  Counter_3_io_reset;
  wire  Counter_3_io_enable;
  wire  _T_1051;
  wire  Counter_4_clock;
  wire  Counter_4_reset;
  wire [63:0] Counter_4_io_out;
  wire  Counter_4_io_reset;
  wire  Counter_4_io_enable;
  wire  SRFF_clock;
  wire  SRFF_reset;
  wire  SRFF_io_input_set;
  wire  SRFF_io_input_reset;
  wire  SRFF_io_input_asyn_reset;
  wire  SRFF_io_output_data;
  wire  _T_1057;
  wire  SRFF_1_clock;
  wire  SRFF_1_reset;
  wire  SRFF_1_io_input_set;
  wire  SRFF_1_io_input_reset;
  wire  SRFF_1_io_input_asyn_reset;
  wire  SRFF_1_io_output_data;
  wire  _T_1064;
  wire  _T_1065;
  reg  _T_1068;
  reg [31:0] _RAND_0;
  wire  _T_1074;
  wire  _T_1075;
  wire  FF_6_clock;
  wire  FF_6_reset;
  wire [31:0] FF_6_io_in;
  wire [31:0] FF_6_io_out;
  wire  FF_6_io_enable;
  wire  _T_1079;
  wire  _T_1080;
  reg  _T_1083;
  reg [31:0] _RAND_1;
  wire  _T_1089;
  wire  _T_1090;
  wire [63:0] _T_1091;
  wire [95:0] _T_1092;
  wire [127:0] _T_1093;
  wire [159:0] _T_1094;
  wire [191:0] _T_1095;
  wire [223:0] _T_1096;
  wire [255:0] _T_1097;
  wire [287:0] _T_1098;
  wire [319:0] _T_1099;
  wire [351:0] _T_1100;
  wire [383:0] _T_1101;
  wire [415:0] _T_1102;
  wire [447:0] _T_1103;
  wire [479:0] _T_1104;
  wire [511:0] _T_1105;
  wire  FF_7_clock;
  wire  FF_7_reset;
  wire [511:0] FF_7_io_in;
  wire [511:0] FF_7_io_out;
  wire  FF_7_io_enable;
  wire  denseStoreBuffers_0_clock;
  wire  denseStoreBuffers_0_reset;
  wire  denseStoreBuffers_0_io_enqVld;
  wire [31:0] denseStoreBuffers_0_io_deq_0;
  wire [31:0] denseStoreBuffers_0_io_deq_1;
  wire [31:0] denseStoreBuffers_0_io_deq_2;
  wire [31:0] denseStoreBuffers_0_io_deq_3;
  wire [31:0] denseStoreBuffers_0_io_deq_4;
  wire [31:0] denseStoreBuffers_0_io_deq_5;
  wire [31:0] denseStoreBuffers_0_io_deq_6;
  wire [31:0] denseStoreBuffers_0_io_deq_7;
  wire [31:0] denseStoreBuffers_0_io_deq_8;
  wire [31:0] denseStoreBuffers_0_io_deq_9;
  wire [31:0] denseStoreBuffers_0_io_deq_10;
  wire [31:0] denseStoreBuffers_0_io_deq_11;
  wire [31:0] denseStoreBuffers_0_io_deq_12;
  wire [31:0] denseStoreBuffers_0_io_deq_13;
  wire [31:0] denseStoreBuffers_0_io_deq_14;
  wire [31:0] denseStoreBuffers_0_io_deq_15;
  wire [63:0] denseStoreBuffers_0_io_deqStrb;
  wire  denseStoreBuffers_0_io_deqVld;
  wire  denseStoreBuffers_0_io_full;
  wire  denseStoreBuffers_0_io_empty;
  wire  denseStoreBuffers_0_io_almostEmpty;
  wire  denseStoreBuffers_0_io_almostFull;
  wire  _T_1109;
  wire  _T_1110;
  wire  _T_1111;
  wire  _T_1112;
  wire  _T_1114;
  wire  _T_1115;
  wire  _T_1116;
  wire  _T_1118;
  wire  _T_1119;
  wire  _T_1120;
  wire  _T_1121;
  wire  _T_1122;
  wire  _T_1123;
  wire  _T_1127;
  wire  _T_1129;
  wire  _T_1130;
  wire  _T_1131;
  wire  _T_1132;
  wire  _T_1133;
  wire  _T_1134;
  wire  _T_1135;
  wire  _T_1136;
  wire  _T_1137;
  wire  _T_1138;
  wire  _T_1139;
  wire  _T_1140;
  wire  _T_1141;
  wire  _T_1142;
  wire  _T_1143;
  wire  _T_1144;
  wire  _T_1145;
  wire  _T_1146;
  wire  _T_1147;
  wire  _T_1148;
  wire  _T_1149;
  wire  _T_1150;
  wire  _T_1151;
  wire  _T_1152;
  wire  _T_1153;
  wire  _T_1154;
  wire  _T_1155;
  wire  _T_1156;
  wire  _T_1157;
  wire  _T_1158;
  wire  _T_1159;
  wire  _T_1160;
  wire  _T_1161;
  wire  _T_1162;
  wire  _T_1163;
  wire  _T_1164;
  wire  _T_1165;
  wire  _T_1166;
  wire  _T_1167;
  wire  _T_1168;
  wire  _T_1169;
  wire  _T_1170;
  wire  _T_1171;
  wire  _T_1172;
  wire  _T_1173;
  wire  _T_1174;
  wire  _T_1175;
  wire  _T_1176;
  wire  _T_1177;
  wire  _T_1178;
  wire  _T_1179;
  wire  _T_1180;
  wire  _T_1181;
  wire  _T_1182;
  wire  _T_1183;
  wire  _T_1184;
  wire  _T_1185;
  wire  _T_1186;
  wire  _T_1187;
  wire  _T_1188;
  wire  _T_1189;
  wire  _T_1190;
  wire  _T_1191;
  wire  _T_1192;
  wire  _T_1193;
  wire  _T_1194;
  wire  Counter_5_clock;
  wire  Counter_5_reset;
  wire [15:0] Counter_5_io_max;
  wire [15:0] Counter_5_io_stride;
  wire [15:0] Counter_5_io_out;
  wire  Counter_5_io_last;
  wire  Counter_5_io_reset;
  wire  Counter_5_io_enable;
  wire  Counter_5_io_done;
  wire  FF_8_clock;
  wire  FF_8_reset;
  wire [15:0] FF_8_io_in;
  wire [15:0] FF_8_io_out;
  wire  FF_8_io_enable;
  wire  _T_1197;
  wire  _T_1202;
  wire  _T_1203;
  wire  FIFOCounter_clock;
  wire  FIFOCounter_reset;
  wire  FIFOCounter_io_enqVld;
  wire  FIFOCounter_io_full;
  wire  FIFOCounter_io_empty;
  wire  _T_1204;
  wire  _T_1205;
  wire  Counter_6_clock;
  wire  Counter_6_reset;
  wire [63:0] Counter_6_io_out;
  wire  Counter_6_io_reset;
  wire  Counter_6_io_enable;
  wire  Counter_7_clock;
  wire  Counter_7_reset;
  wire [63:0] Counter_7_io_out;
  wire  Counter_7_io_reset;
  wire  Counter_7_io_enable;
  wire  Counter_8_clock;
  wire  Counter_8_reset;
  wire [63:0] Counter_8_io_out;
  wire  Counter_8_io_reset;
  wire  Counter_8_io_enable;
  wire  burstCounterMaxLatch_clock;
  wire  burstCounterMaxLatch_reset;
  wire [31:0] burstCounterMaxLatch_io_in;
  wire [31:0] burstCounterMaxLatch_io_out;
  wire  burstCounterMaxLatch_io_enable;
  wire [31:0] burstCounterMax;
  wire  _T_1227;
  wire  _T_1229;
  wire [31:0] _T_1231;
  wire  _T_1233;
  wire  _T_1235;
  wire  dramReadyFF_clock;
  wire  dramReadyFF_reset;
  wire  dramReadyFF_io_in;
  wire  dramReadyFF_io_init;
  wire  dramReadyFF_io_reset;
  wire  dramReadyFF_io_out;
  wire  dramReadyFF_io_enable;
  wire  dramReadyFFEnabler;
  wire  _T_1243;
  wire  _T_1244;
  wire  _T_1246;
  wire  _T_1247;
  wire  _T_1249;
  wire  _T_1255;
  wire  _T_1256;
  wire  cycleCount_clock;
  wire  cycleCount_reset;
  wire [63:0] cycleCount_io_out;
  wire  cycleCount_io_reset;
  wire  cycleCount_io_enable;
  wire  _T_1261;
  wire  rdataEnqCount_clock;
  wire  rdataEnqCount_reset;
  wire [63:0] rdataEnqCount_io_out;
  wire  rdataEnqCount_io_reset;
  wire  rdataEnqCount_io_enable;
  wire  _T_1266;
  wire  _T_1267;
  wire  wdataCount_clock;
  wire  wdataCount_reset;
  wire [63:0] wdataCount_io_out;
  wire  wdataCount_io_reset;
  wire  wdataCount_io_enable;
  wire  _T_1272;
  wire  _T_1273;
  wire  Counter_9_clock;
  wire  Counter_9_reset;
  wire [63:0] Counter_9_io_out;
  wire  Counter_9_io_reset;
  wire  Counter_9_io_enable;
  wire  _T_1278;
  wire  _T_1279;
  wire  _T_1280;
  wire  _T_1281;
  wire  _T_1282;
  wire  Counter_10_clock;
  wire  Counter_10_reset;
  wire [63:0] Counter_10_io_out;
  wire  Counter_10_io_reset;
  wire  Counter_10_io_enable;
  wire  _T_1290;
  wire  Counter_11_clock;
  wire  Counter_11_reset;
  wire [63:0] Counter_11_io_out;
  wire  Counter_11_io_reset;
  wire  Counter_11_io_enable;
  wire  _T_1295;
  wire  Counter_12_clock;
  wire  Counter_12_reset;
  wire [63:0] Counter_12_io_out;
  wire  Counter_12_io_reset;
  wire  Counter_12_io_enable;
  wire  _T_1301;
  wire  Counter_13_clock;
  wire  Counter_13_reset;
  wire [63:0] Counter_13_io_out;
  wire  Counter_13_io_reset;
  wire  Counter_13_io_enable;
  wire  _T_1308;
  wire  _T_1309;
  wire  Counter_14_clock;
  wire  Counter_14_reset;
  wire [63:0] Counter_14_io_out;
  wire  Counter_14_io_reset;
  wire  Counter_14_io_enable;
  wire  _T_1316;
  wire  Counter_15_clock;
  wire  Counter_15_reset;
  wire [63:0] Counter_15_io_out;
  wire  Counter_15_io_reset;
  wire  Counter_15_io_enable;
  wire  Counter_16_clock;
  wire  Counter_16_reset;
  wire [63:0] Counter_16_io_out;
  wire  Counter_16_io_reset;
  wire  Counter_16_io_enable;
  wire  Counter_17_clock;
  wire  Counter_17_reset;
  wire [63:0] Counter_17_io_out;
  wire  Counter_17_io_reset;
  wire  Counter_17_io_enable;
  wire  _T_1335;
  wire  Counter_18_clock;
  wire  Counter_18_reset;
  wire [63:0] Counter_18_io_out;
  wire  Counter_18_io_reset;
  wire  Counter_18_io_enable;
  wire  Counter_19_clock;
  wire  Counter_19_reset;
  wire [63:0] Counter_19_io_out;
  wire  Counter_19_io_reset;
  wire  Counter_19_io_enable;
  wire  _T_1345;
  wire  _T_1346;
  wire  _T_1347;
  wire  Counter_20_clock;
  wire  Counter_20_reset;
  wire [63:0] Counter_20_io_out;
  wire  Counter_20_io_reset;
  wire  Counter_20_io_enable;
  wire  _T_1352;
  wire  _T_1353;
  wire  _T_1354;
  wire  Counter_21_clock;
  wire  Counter_21_reset;
  wire [63:0] Counter_21_io_out;
  wire  Counter_21_io_reset;
  wire  Counter_21_io_enable;
  wire  _T_1362;
  wire  Counter_22_clock;
  wire  Counter_22_reset;
  wire [63:0] Counter_22_io_out;
  wire  Counter_22_io_reset;
  wire  Counter_22_io_enable;
  wire  _T_1367;
  wire  Counter_23_clock;
  wire  Counter_23_reset;
  wire [63:0] Counter_23_io_out;
  wire  Counter_23_io_reset;
  wire  Counter_23_io_enable;
  wire  _T_1372;
  wire  _T_1373;
  wire  _T_1374;
  wire  Counter_24_clock;
  wire  Counter_24_reset;
  wire [63:0] Counter_24_io_out;
  wire  Counter_24_io_reset;
  wire  Counter_24_io_enable;
  wire  _T_1379;
  wire  _T_1380;
  wire  _T_1381;
  wire  Counter_25_clock;
  wire  Counter_25_reset;
  wire [63:0] Counter_25_io_out;
  wire  Counter_25_io_reset;
  wire  Counter_25_io_enable;
  wire  _T_1389;
  wire  Counter_26_clock;
  wire  Counter_26_reset;
  wire [63:0] Counter_26_io_out;
  wire  Counter_26_io_reset;
  wire  Counter_26_io_enable;
  wire  Counter_27_clock;
  wire  Counter_27_reset;
  wire [63:0] Counter_27_io_out;
  wire  Counter_27_io_reset;
  wire  Counter_27_io_enable;
  wire  Counter_28_clock;
  wire  Counter_28_reset;
  wire [63:0] Counter_28_io_out;
  wire  Counter_28_io_reset;
  wire  Counter_28_io_enable;
  wire  Counter_29_clock;
  wire  Counter_29_reset;
  wire [63:0] Counter_29_io_out;
  wire  Counter_29_io_reset;
  wire  Counter_29_io_enable;
  wire  Counter_30_clock;
  wire  Counter_30_reset;
  wire [63:0] Counter_30_io_out;
  wire  Counter_30_io_reset;
  wire  Counter_30_io_enable;
  wire  Counter_31_clock;
  wire  Counter_31_reset;
  wire [63:0] Counter_31_io_out;
  wire  Counter_31_io_reset;
  wire  Counter_31_io_enable;
  wire  Counter_32_clock;
  wire  Counter_32_reset;
  wire [63:0] Counter_32_io_out;
  wire  Counter_32_io_reset;
  wire  Counter_32_io_enable;
  wire  Counter_33_clock;
  wire  Counter_33_reset;
  wire [63:0] Counter_33_io_out;
  wire  Counter_33_io_reset;
  wire  Counter_33_io_enable;
  wire  _T_1425;
  wire  Counter_34_clock;
  wire  Counter_34_reset;
  wire [63:0] Counter_34_io_out;
  wire  Counter_34_io_reset;
  wire  Counter_34_io_enable;
  wire  FF_9_clock;
  wire  FF_9_reset;
  wire [5:0] FF_9_io_in;
  wire [5:0] FF_9_io_out;
  wire  FF_9_io_enable;
  wire  Counter_35_clock;
  wire  Counter_35_reset;
  wire [63:0] Counter_35_io_out;
  wire  Counter_35_io_reset;
  wire  Counter_35_io_enable;
  wire  Counter_36_clock;
  wire  Counter_36_reset;
  wire [63:0] Counter_36_io_out;
  wire  Counter_36_io_reset;
  wire  Counter_36_io_enable;
  wire  _T_1443;
  wire  Counter_37_clock;
  wire  Counter_37_reset;
  wire [63:0] Counter_37_io_out;
  wire  Counter_37_io_reset;
  wire  Counter_37_io_enable;
  wire  _T_1448;
  wire  Counter_38_clock;
  wire  Counter_38_reset;
  wire [63:0] Counter_38_io_out;
  wire  Counter_38_io_reset;
  wire  Counter_38_io_enable;
  wire  Counter_39_clock;
  wire  Counter_39_reset;
  wire [63:0] Counter_39_io_out;
  wire  Counter_39_io_reset;
  wire  Counter_39_io_enable;
  wire  Counter_40_clock;
  wire  Counter_40_reset;
  wire [63:0] Counter_40_io_out;
  wire  Counter_40_io_reset;
  wire  Counter_40_io_enable;
  wire  Counter_41_clock;
  wire  Counter_41_reset;
  wire [63:0] Counter_41_io_out;
  wire  Counter_41_io_reset;
  wire  Counter_41_io_enable;
  wire  Counter_42_clock;
  wire  Counter_42_reset;
  wire [63:0] Counter_42_io_out;
  wire  Counter_42_io_reset;
  wire  Counter_42_io_enable;
  wire  _T_1469;
  wire  Counter_43_clock;
  wire  Counter_43_reset;
  wire [63:0] Counter_43_io_out;
  wire  Counter_43_io_reset;
  wire  Counter_43_io_enable;
  wire  Counter_44_clock;
  wire  Counter_44_reset;
  wire [63:0] Counter_44_io_out;
  wire  Counter_44_io_reset;
  wire  Counter_44_io_enable;
  wire  _T_1480;
  wire  Counter_45_clock;
  wire  Counter_45_reset;
  wire [63:0] Counter_45_io_out;
  wire  Counter_45_io_reset;
  wire  Counter_45_io_enable;
  wire  _T_1486;
  wire  Counter_46_clock;
  wire  Counter_46_reset;
  wire [63:0] Counter_46_io_out;
  wire  Counter_46_io_reset;
  wire  Counter_46_io_enable;
  wire  Counter_47_clock;
  wire  Counter_47_reset;
  wire [63:0] Counter_47_io_out;
  wire  Counter_47_io_reset;
  wire  Counter_47_io_enable;
  wire  Counter_48_clock;
  wire  Counter_48_reset;
  wire [63:0] Counter_48_io_out;
  wire  Counter_48_io_reset;
  wire  Counter_48_io_enable;
  wire  Counter_49_clock;
  wire  Counter_49_reset;
  wire [63:0] Counter_49_io_out;
  wire  Counter_49_io_reset;
  wire  Counter_49_io_enable;
  wire  Counter_50_clock;
  wire  Counter_50_reset;
  wire [63:0] Counter_50_io_out;
  wire  Counter_50_io_reset;
  wire  Counter_50_io_enable;
  wire  Counter_51_clock;
  wire  Counter_51_reset;
  wire [63:0] Counter_51_io_out;
  wire  Counter_51_io_reset;
  wire  Counter_51_io_enable;
  wire  Counter_52_clock;
  wire  Counter_52_reset;
  wire [63:0] Counter_52_io_out;
  wire  Counter_52_io_reset;
  wire  Counter_52_io_enable;
  wire  Counter_53_clock;
  wire  Counter_53_reset;
  wire [63:0] Counter_53_io_out;
  wire  Counter_53_io_reset;
  wire  Counter_53_io_enable;
  wire  Counter_54_clock;
  wire  Counter_54_reset;
  wire [63:0] Counter_54_io_out;
  wire  Counter_54_io_reset;
  wire  Counter_54_io_enable;
  wire  Counter_55_clock;
  wire  Counter_55_reset;
  wire [63:0] Counter_55_io_out;
  wire  Counter_55_io_reset;
  wire  Counter_55_io_enable;
  wire  Counter_56_clock;
  wire  Counter_56_reset;
  wire [63:0] Counter_56_io_out;
  wire  Counter_56_io_reset;
  wire  Counter_56_io_enable;
  wire  Counter_57_clock;
  wire  Counter_57_reset;
  wire [63:0] Counter_57_io_out;
  wire  Counter_57_io_reset;
  wire  Counter_57_io_enable;
  wire  Counter_58_clock;
  wire  Counter_58_reset;
  wire [63:0] Counter_58_io_out;
  wire  Counter_58_io_reset;
  wire  Counter_58_io_enable;
  wire  Counter_59_clock;
  wire  Counter_59_reset;
  wire [63:0] Counter_59_io_out;
  wire  Counter_59_io_reset;
  wire  Counter_59_io_enable;
  wire  FF_10_clock;
  wire  FF_10_reset;
  wire [63:0] FF_10_io_in;
  wire [63:0] FF_10_io_init;
  wire  FF_10_io_reset;
  wire [63:0] FF_10_io_out;
  wire  FF_10_io_enable;
  wire  FF_11_clock;
  wire  FF_11_reset;
  wire [7:0] FF_11_io_in;
  wire [7:0] FF_11_io_out;
  wire  FF_11_io_enable;
  wire  FF_12_clock;
  wire  FF_12_reset;
  wire [2:0] FF_12_io_in;
  wire [2:0] FF_12_io_out;
  wire  FF_12_io_enable;
  wire  FF_13_clock;
  wire  FF_13_reset;
  wire  FF_13_io_in;
  wire  FF_13_io_init;
  wire  FF_13_io_reset;
  wire  FF_13_io_out;
  wire  FF_13_io_enable;
  wire  FF_14_clock;
  wire  FF_14_reset;
  wire [1:0] FF_14_io_in;
  wire [1:0] FF_14_io_out;
  wire  FF_14_io_enable;
  wire  FF_15_clock;
  wire  FF_15_reset;
  wire [63:0] FF_15_io_in;
  wire [63:0] FF_15_io_init;
  wire  FF_15_io_reset;
  wire [63:0] FF_15_io_out;
  wire  FF_15_io_enable;
  wire  FF_16_clock;
  wire  FF_16_reset;
  wire [7:0] FF_16_io_in;
  wire [7:0] FF_16_io_out;
  wire  FF_16_io_enable;
  wire  FF_17_clock;
  wire  FF_17_reset;
  wire [511:0] FF_17_io_in;
  wire [511:0] FF_17_io_out;
  wire  FF_17_io_enable;
  wire  FF_18_clock;
  wire  FF_18_reset;
  wire [63:0] FF_18_io_in;
  wire [63:0] FF_18_io_init;
  wire  FF_18_io_reset;
  wire [63:0] FF_18_io_out;
  wire  FF_18_io_enable;
  wire  FF_19_clock;
  wire  FF_19_reset;
  wire [511:0] FF_19_io_in;
  wire [511:0] FF_19_io_out;
  wire  FF_19_io_enable;
  wire  FF_20_clock;
  wire  FF_20_reset;
  wire [63:0] FF_20_io_in;
  wire [63:0] FF_20_io_init;
  wire  FF_20_io_reset;
  wire [63:0] FF_20_io_out;
  wire  FF_20_io_enable;
  wire  FF_21_clock;
  wire  FF_21_reset;
  wire [511:0] FF_21_io_in;
  wire [511:0] FF_21_io_out;
  wire  FF_21_io_enable;
  wire  FF_22_clock;
  wire  FF_22_reset;
  wire [63:0] FF_22_io_in;
  wire [63:0] FF_22_io_init;
  wire  FF_22_io_reset;
  wire [63:0] FF_22_io_out;
  wire  FF_22_io_enable;
  wire  Counter_60_clock;
  wire  Counter_60_reset;
  wire [63:0] Counter_60_io_out;
  wire  Counter_60_io_reset;
  wire  Counter_60_io_enable;
  wire  Counter_61_clock;
  wire  Counter_61_reset;
  wire [63:0] Counter_61_io_out;
  wire  Counter_61_io_reset;
  wire  Counter_61_io_enable;
  wire  Counter_62_clock;
  wire  Counter_62_reset;
  wire [63:0] Counter_62_io_out;
  wire  Counter_62_io_reset;
  wire  Counter_62_io_enable;
  wire  Counter_63_clock;
  wire  Counter_63_reset;
  wire [63:0] Counter_63_io_out;
  wire  Counter_63_io_reset;
  wire  Counter_63_io_enable;
  wire  Counter_64_clock;
  wire  Counter_64_reset;
  wire [63:0] Counter_64_io_out;
  wire  Counter_64_io_reset;
  wire  Counter_64_io_enable;
  wire  Counter_65_clock;
  wire  Counter_65_reset;
  wire [63:0] Counter_65_io_out;
  wire  Counter_65_io_reset;
  wire  Counter_65_io_enable;
  wire  Counter_66_clock;
  wire  Counter_66_reset;
  wire [63:0] Counter_66_io_out;
  wire  Counter_66_io_reset;
  wire  Counter_66_io_enable;
  wire  Counter_67_clock;
  wire  Counter_67_reset;
  wire [63:0] Counter_67_io_out;
  wire  Counter_67_io_reset;
  wire  Counter_67_io_enable;
  wire  Counter_68_clock;
  wire  Counter_68_reset;
  wire [63:0] Counter_68_io_out;
  wire  Counter_68_io_reset;
  wire  Counter_68_io_enable;
  wire  Counter_69_clock;
  wire  Counter_69_reset;
  wire [63:0] Counter_69_io_out;
  wire  Counter_69_io_reset;
  wire  Counter_69_io_enable;
  wire  Counter_70_clock;
  wire  Counter_70_reset;
  wire [63:0] Counter_70_io_out;
  wire  Counter_70_io_reset;
  wire  Counter_70_io_enable;
  wire  Counter_71_clock;
  wire  Counter_71_reset;
  wire [63:0] Counter_71_io_out;
  wire  Counter_71_io_reset;
  wire  Counter_71_io_enable;
  wire  Counter_72_clock;
  wire  Counter_72_reset;
  wire [63:0] Counter_72_io_out;
  wire  Counter_72_io_reset;
  wire  Counter_72_io_enable;
  wire  FF_23_clock;
  wire  FF_23_reset;
  wire [63:0] FF_23_io_in;
  wire [63:0] FF_23_io_init;
  wire  FF_23_io_reset;
  wire [63:0] FF_23_io_out;
  wire  FF_23_io_enable;
  wire  FF_24_clock;
  wire  FF_24_reset;
  wire [7:0] FF_24_io_in;
  wire [7:0] FF_24_io_out;
  wire  FF_24_io_enable;
  wire  FF_25_clock;
  wire  FF_25_reset;
  wire [2:0] FF_25_io_in;
  wire [2:0] FF_25_io_out;
  wire  FF_25_io_enable;
  wire  FF_26_clock;
  wire  FF_26_reset;
  wire [1:0] FF_26_io_in;
  wire [1:0] FF_26_io_out;
  wire  FF_26_io_enable;
  wire  FF_27_clock;
  wire  FF_27_reset;
  wire [63:0] FF_27_io_in;
  wire [63:0] FF_27_io_init;
  wire  FF_27_io_reset;
  wire [63:0] FF_27_io_out;
  wire  FF_27_io_enable;
  wire  FF_28_clock;
  wire  FF_28_reset;
  wire [7:0] FF_28_io_in;
  wire [7:0] FF_28_io_out;
  wire  FF_28_io_enable;
  wire  FF_29_clock;
  wire  FF_29_reset;
  wire [511:0] FF_29_io_in;
  wire [511:0] FF_29_io_out;
  wire  FF_29_io_enable;
  wire  FF_30_clock;
  wire  FF_30_reset;
  wire [63:0] FF_30_io_in;
  wire [63:0] FF_30_io_init;
  wire  FF_30_io_reset;
  wire [63:0] FF_30_io_out;
  wire  FF_30_io_enable;
  wire  FF_31_clock;
  wire  FF_31_reset;
  wire [511:0] FF_31_io_in;
  wire [511:0] FF_31_io_out;
  wire  FF_31_io_enable;
  wire  FF_32_clock;
  wire  FF_32_reset;
  wire [63:0] FF_32_io_in;
  wire [63:0] FF_32_io_init;
  wire  FF_32_io_reset;
  wire [63:0] FF_32_io_out;
  wire  FF_32_io_enable;
  wire  FF_33_clock;
  wire  FF_33_reset;
  wire [511:0] FF_33_io_in;
  wire [511:0] FF_33_io_out;
  wire  FF_33_io_enable;
  wire  FF_34_clock;
  wire  FF_34_reset;
  wire [63:0] FF_34_io_in;
  wire [63:0] FF_34_io_init;
  wire  FF_34_io_reset;
  wire [63:0] FF_34_io_out;
  wire  FF_34_io_enable;
  FIFOArbiter cmdArbiter (
    .clock(cmdArbiter_clock),
    .reset(cmdArbiter_reset),
    .io_fifo_0_enq_0_addr(cmdArbiter_io_fifo_0_enq_0_addr),
    .io_fifo_0_enq_0_isWr(cmdArbiter_io_fifo_0_enq_0_isWr),
    .io_fifo_0_enq_0_size(cmdArbiter_io_fifo_0_enq_0_size),
    .io_fifo_0_enqVld(cmdArbiter_io_fifo_0_enqVld),
    .io_fifo_0_deq_0_addr(cmdArbiter_io_fifo_0_deq_0_addr),
    .io_fifo_0_deq_0_isWr(cmdArbiter_io_fifo_0_deq_0_isWr),
    .io_fifo_0_deq_0_size(cmdArbiter_io_fifo_0_deq_0_size),
    .io_fifo_0_deqVld(cmdArbiter_io_fifo_0_deqVld),
    .io_fifo_0_full(cmdArbiter_io_fifo_0_full),
    .io_fifo_0_empty(cmdArbiter_io_fifo_0_empty),
    .io_fifo_0_almostEmpty(cmdArbiter_io_fifo_0_almostEmpty),
    .io_fifo_1_deq_0_addr(cmdArbiter_io_fifo_1_deq_0_addr),
    .io_fifo_1_deq_0_isWr(cmdArbiter_io_fifo_1_deq_0_isWr),
    .io_fifo_1_deq_0_size(cmdArbiter_io_fifo_1_deq_0_size),
    .io_fifo_1_deqVld(cmdArbiter_io_fifo_1_deqVld),
    .io_fifo_1_empty(cmdArbiter_io_fifo_1_empty),
    .io_enq_0_0_addr(cmdArbiter_io_enq_0_0_addr),
    .io_enq_0_0_isWr(cmdArbiter_io_enq_0_0_isWr),
    .io_enq_0_0_size(cmdArbiter_io_enq_0_0_size),
    .io_enqVld_0(cmdArbiter_io_enqVld_0),
    .io_full_0(cmdArbiter_io_full_0),
    .io_deq_0_addr(cmdArbiter_io_deq_0_addr),
    .io_deq_0_isWr(cmdArbiter_io_deq_0_isWr),
    .io_deq_0_size(cmdArbiter_io_deq_0_size),
    .io_deqVld(cmdArbiter_io_deqVld),
    .io_deqReady(cmdArbiter_io_deqReady),
    .io_empty(cmdArbiter_io_empty),
    .io_tag(cmdArbiter_io_tag)
  );
  FIFOCore cmdFifos_0 (
    .clock(cmdFifos_0_clock),
    .reset(cmdFifos_0_reset),
    .io_enq_0_addr(cmdFifos_0_io_enq_0_addr),
    .io_enq_0_isWr(cmdFifos_0_io_enq_0_isWr),
    .io_enq_0_size(cmdFifos_0_io_enq_0_size),
    .io_enqVld(cmdFifos_0_io_enqVld),
    .io_deq_0_addr(cmdFifos_0_io_deq_0_addr),
    .io_deq_0_isWr(cmdFifos_0_io_deq_0_isWr),
    .io_deq_0_size(cmdFifos_0_io_deq_0_size),
    .io_deqVld(cmdFifos_0_io_deqVld),
    .io_full(cmdFifos_0_io_full),
    .io_empty(cmdFifos_0_io_empty),
    .io_almostEmpty(cmdFifos_0_io_almostEmpty)
  );
  FIFOCore cmdFifos_1 (
    .clock(cmdFifos_1_clock),
    .reset(cmdFifos_1_reset),
    .io_enq_0_addr(cmdFifos_1_io_enq_0_addr),
    .io_enq_0_isWr(cmdFifos_1_io_enq_0_isWr),
    .io_enq_0_size(cmdFifos_1_io_enq_0_size),
    .io_enqVld(cmdFifos_1_io_enqVld),
    .io_deq_0_addr(cmdFifos_1_io_deq_0_addr),
    .io_deq_0_isWr(cmdFifos_1_io_deq_0_isWr),
    .io_deq_0_size(cmdFifos_1_io_deq_0_size),
    .io_deqVld(cmdFifos_1_io_deqVld),
    .io_full(cmdFifos_1_io_full),
    .io_empty(cmdFifos_1_io_empty),
    .io_almostEmpty(cmdFifos_1_io_almostEmpty)
  );
  FF_136 FF (
    .clock(FF_clock),
    .reset(FF_reset),
    .io_in(FF_io_in),
    .io_init(FF_io_init),
    .io_reset(FF_io_reset),
    .io_out(FF_io_out),
    .io_enable(FF_io_enable)
  );
  Counter_15 sizeCounter (
    .clock(sizeCounter_clock),
    .reset(sizeCounter_reset),
    .io_max(sizeCounter_io_max),
    .io_stride(sizeCounter_io_stride),
    .io_out(sizeCounter_io_out),
    .io_last(sizeCounter_io_last),
    .io_reset(sizeCounter_io_reset),
    .io_enable(sizeCounter_io_enable),
    .io_done(sizeCounter_io_done)
  );
  MuxN_4 isSparseMux (
    .io_ins_0(isSparseMux_io_ins_0),
    .io_ins_1(isSparseMux_io_ins_1),
    .io_sel(isSparseMux_io_sel),
    .io_out(isSparseMux_io_out)
  );
  Counter_15 burstCounter (
    .clock(burstCounter_clock),
    .reset(burstCounter_reset),
    .io_max(burstCounter_io_max),
    .io_stride(burstCounter_io_stride),
    .io_out(burstCounter_io_out),
    .io_last(burstCounter_io_last),
    .io_reset(burstCounter_io_reset),
    .io_enable(burstCounter_io_enable),
    .io_done(burstCounter_io_done)
  );
  Counter_17 burstTagCounter (
    .clock(burstTagCounter_clock),
    .reset(burstTagCounter_reset),
    .io_out(burstTagCounter_io_out),
    .io_reset(burstTagCounter_io_reset),
    .io_enable(burstTagCounter_io_enable)
  );
  FF_115 cmdCooldown (
    .clock(cmdCooldown_clock),
    .reset(cmdCooldown_reset),
    .io_in(cmdCooldown_io_in),
    .io_init(cmdCooldown_io_init),
    .io_reset(cmdCooldown_io_reset),
    .io_out(cmdCooldown_io_out),
    .io_enable(cmdCooldown_io_enable)
  );
  FF_115 burstCounterDoneLatch (
    .clock(burstCounterDoneLatch_clock),
    .reset(burstCounterDoneLatch_reset),
    .io_in(burstCounterDoneLatch_io_in),
    .io_init(burstCounterDoneLatch_io_init),
    .io_reset(burstCounterDoneLatch_io_reset),
    .io_out(burstCounterDoneLatch_io_out),
    .io_enable(burstCounterDoneLatch_io_enable)
  );
  FF_115 sizeCounterDoneLatch (
    .clock(sizeCounterDoneLatch_clock),
    .reset(sizeCounterDoneLatch_reset),
    .io_in(sizeCounterDoneLatch_io_in),
    .io_init(sizeCounterDoneLatch_io_init),
    .io_reset(sizeCounterDoneLatch_io_reset),
    .io_out(sizeCounterDoneLatch_io_out),
    .io_enable(sizeCounterDoneLatch_io_enable)
  );
  MuxN_5 rrespReadyMux (
    .io_ins_0(rrespReadyMux_io_ins_0),
    .io_out(rrespReadyMux_io_out)
  );
  MuxN_6 wdataMux (
    .io_ins_0_valid(wdataMux_io_ins_0_valid),
    .io_ins_0_bits_wdata_0(wdataMux_io_ins_0_bits_wdata_0),
    .io_ins_0_bits_wdata_1(wdataMux_io_ins_0_bits_wdata_1),
    .io_ins_0_bits_wdata_2(wdataMux_io_ins_0_bits_wdata_2),
    .io_ins_0_bits_wdata_3(wdataMux_io_ins_0_bits_wdata_3),
    .io_ins_0_bits_wdata_4(wdataMux_io_ins_0_bits_wdata_4),
    .io_ins_0_bits_wdata_5(wdataMux_io_ins_0_bits_wdata_5),
    .io_ins_0_bits_wdata_6(wdataMux_io_ins_0_bits_wdata_6),
    .io_ins_0_bits_wdata_7(wdataMux_io_ins_0_bits_wdata_7),
    .io_ins_0_bits_wdata_8(wdataMux_io_ins_0_bits_wdata_8),
    .io_ins_0_bits_wdata_9(wdataMux_io_ins_0_bits_wdata_9),
    .io_ins_0_bits_wdata_10(wdataMux_io_ins_0_bits_wdata_10),
    .io_ins_0_bits_wdata_11(wdataMux_io_ins_0_bits_wdata_11),
    .io_ins_0_bits_wdata_12(wdataMux_io_ins_0_bits_wdata_12),
    .io_ins_0_bits_wdata_13(wdataMux_io_ins_0_bits_wdata_13),
    .io_ins_0_bits_wdata_14(wdataMux_io_ins_0_bits_wdata_14),
    .io_ins_0_bits_wdata_15(wdataMux_io_ins_0_bits_wdata_15),
    .io_ins_0_bits_wstrb_0(wdataMux_io_ins_0_bits_wstrb_0),
    .io_ins_0_bits_wstrb_1(wdataMux_io_ins_0_bits_wstrb_1),
    .io_ins_0_bits_wstrb_2(wdataMux_io_ins_0_bits_wstrb_2),
    .io_ins_0_bits_wstrb_3(wdataMux_io_ins_0_bits_wstrb_3),
    .io_ins_0_bits_wstrb_4(wdataMux_io_ins_0_bits_wstrb_4),
    .io_ins_0_bits_wstrb_5(wdataMux_io_ins_0_bits_wstrb_5),
    .io_ins_0_bits_wstrb_6(wdataMux_io_ins_0_bits_wstrb_6),
    .io_ins_0_bits_wstrb_7(wdataMux_io_ins_0_bits_wstrb_7),
    .io_ins_0_bits_wstrb_8(wdataMux_io_ins_0_bits_wstrb_8),
    .io_ins_0_bits_wstrb_9(wdataMux_io_ins_0_bits_wstrb_9),
    .io_ins_0_bits_wstrb_10(wdataMux_io_ins_0_bits_wstrb_10),
    .io_ins_0_bits_wstrb_11(wdataMux_io_ins_0_bits_wstrb_11),
    .io_ins_0_bits_wstrb_12(wdataMux_io_ins_0_bits_wstrb_12),
    .io_ins_0_bits_wstrb_13(wdataMux_io_ins_0_bits_wstrb_13),
    .io_ins_0_bits_wstrb_14(wdataMux_io_ins_0_bits_wstrb_14),
    .io_ins_0_bits_wstrb_15(wdataMux_io_ins_0_bits_wstrb_15),
    .io_ins_0_bits_wstrb_16(wdataMux_io_ins_0_bits_wstrb_16),
    .io_ins_0_bits_wstrb_17(wdataMux_io_ins_0_bits_wstrb_17),
    .io_ins_0_bits_wstrb_18(wdataMux_io_ins_0_bits_wstrb_18),
    .io_ins_0_bits_wstrb_19(wdataMux_io_ins_0_bits_wstrb_19),
    .io_ins_0_bits_wstrb_20(wdataMux_io_ins_0_bits_wstrb_20),
    .io_ins_0_bits_wstrb_21(wdataMux_io_ins_0_bits_wstrb_21),
    .io_ins_0_bits_wstrb_22(wdataMux_io_ins_0_bits_wstrb_22),
    .io_ins_0_bits_wstrb_23(wdataMux_io_ins_0_bits_wstrb_23),
    .io_ins_0_bits_wstrb_24(wdataMux_io_ins_0_bits_wstrb_24),
    .io_ins_0_bits_wstrb_25(wdataMux_io_ins_0_bits_wstrb_25),
    .io_ins_0_bits_wstrb_26(wdataMux_io_ins_0_bits_wstrb_26),
    .io_ins_0_bits_wstrb_27(wdataMux_io_ins_0_bits_wstrb_27),
    .io_ins_0_bits_wstrb_28(wdataMux_io_ins_0_bits_wstrb_28),
    .io_ins_0_bits_wstrb_29(wdataMux_io_ins_0_bits_wstrb_29),
    .io_ins_0_bits_wstrb_30(wdataMux_io_ins_0_bits_wstrb_30),
    .io_ins_0_bits_wstrb_31(wdataMux_io_ins_0_bits_wstrb_31),
    .io_ins_0_bits_wstrb_32(wdataMux_io_ins_0_bits_wstrb_32),
    .io_ins_0_bits_wstrb_33(wdataMux_io_ins_0_bits_wstrb_33),
    .io_ins_0_bits_wstrb_34(wdataMux_io_ins_0_bits_wstrb_34),
    .io_ins_0_bits_wstrb_35(wdataMux_io_ins_0_bits_wstrb_35),
    .io_ins_0_bits_wstrb_36(wdataMux_io_ins_0_bits_wstrb_36),
    .io_ins_0_bits_wstrb_37(wdataMux_io_ins_0_bits_wstrb_37),
    .io_ins_0_bits_wstrb_38(wdataMux_io_ins_0_bits_wstrb_38),
    .io_ins_0_bits_wstrb_39(wdataMux_io_ins_0_bits_wstrb_39),
    .io_ins_0_bits_wstrb_40(wdataMux_io_ins_0_bits_wstrb_40),
    .io_ins_0_bits_wstrb_41(wdataMux_io_ins_0_bits_wstrb_41),
    .io_ins_0_bits_wstrb_42(wdataMux_io_ins_0_bits_wstrb_42),
    .io_ins_0_bits_wstrb_43(wdataMux_io_ins_0_bits_wstrb_43),
    .io_ins_0_bits_wstrb_44(wdataMux_io_ins_0_bits_wstrb_44),
    .io_ins_0_bits_wstrb_45(wdataMux_io_ins_0_bits_wstrb_45),
    .io_ins_0_bits_wstrb_46(wdataMux_io_ins_0_bits_wstrb_46),
    .io_ins_0_bits_wstrb_47(wdataMux_io_ins_0_bits_wstrb_47),
    .io_ins_0_bits_wstrb_48(wdataMux_io_ins_0_bits_wstrb_48),
    .io_ins_0_bits_wstrb_49(wdataMux_io_ins_0_bits_wstrb_49),
    .io_ins_0_bits_wstrb_50(wdataMux_io_ins_0_bits_wstrb_50),
    .io_ins_0_bits_wstrb_51(wdataMux_io_ins_0_bits_wstrb_51),
    .io_ins_0_bits_wstrb_52(wdataMux_io_ins_0_bits_wstrb_52),
    .io_ins_0_bits_wstrb_53(wdataMux_io_ins_0_bits_wstrb_53),
    .io_ins_0_bits_wstrb_54(wdataMux_io_ins_0_bits_wstrb_54),
    .io_ins_0_bits_wstrb_55(wdataMux_io_ins_0_bits_wstrb_55),
    .io_ins_0_bits_wstrb_56(wdataMux_io_ins_0_bits_wstrb_56),
    .io_ins_0_bits_wstrb_57(wdataMux_io_ins_0_bits_wstrb_57),
    .io_ins_0_bits_wstrb_58(wdataMux_io_ins_0_bits_wstrb_58),
    .io_ins_0_bits_wstrb_59(wdataMux_io_ins_0_bits_wstrb_59),
    .io_ins_0_bits_wstrb_60(wdataMux_io_ins_0_bits_wstrb_60),
    .io_ins_0_bits_wstrb_61(wdataMux_io_ins_0_bits_wstrb_61),
    .io_ins_0_bits_wstrb_62(wdataMux_io_ins_0_bits_wstrb_62),
    .io_ins_0_bits_wstrb_63(wdataMux_io_ins_0_bits_wstrb_63),
    .io_out_valid(wdataMux_io_out_valid),
    .io_out_bits_wdata_0(wdataMux_io_out_bits_wdata_0),
    .io_out_bits_wdata_1(wdataMux_io_out_bits_wdata_1),
    .io_out_bits_wdata_2(wdataMux_io_out_bits_wdata_2),
    .io_out_bits_wdata_3(wdataMux_io_out_bits_wdata_3),
    .io_out_bits_wdata_4(wdataMux_io_out_bits_wdata_4),
    .io_out_bits_wdata_5(wdataMux_io_out_bits_wdata_5),
    .io_out_bits_wdata_6(wdataMux_io_out_bits_wdata_6),
    .io_out_bits_wdata_7(wdataMux_io_out_bits_wdata_7),
    .io_out_bits_wdata_8(wdataMux_io_out_bits_wdata_8),
    .io_out_bits_wdata_9(wdataMux_io_out_bits_wdata_9),
    .io_out_bits_wdata_10(wdataMux_io_out_bits_wdata_10),
    .io_out_bits_wdata_11(wdataMux_io_out_bits_wdata_11),
    .io_out_bits_wdata_12(wdataMux_io_out_bits_wdata_12),
    .io_out_bits_wdata_13(wdataMux_io_out_bits_wdata_13),
    .io_out_bits_wdata_14(wdataMux_io_out_bits_wdata_14),
    .io_out_bits_wdata_15(wdataMux_io_out_bits_wdata_15),
    .io_out_bits_wstrb_0(wdataMux_io_out_bits_wstrb_0),
    .io_out_bits_wstrb_1(wdataMux_io_out_bits_wstrb_1),
    .io_out_bits_wstrb_2(wdataMux_io_out_bits_wstrb_2),
    .io_out_bits_wstrb_3(wdataMux_io_out_bits_wstrb_3),
    .io_out_bits_wstrb_4(wdataMux_io_out_bits_wstrb_4),
    .io_out_bits_wstrb_5(wdataMux_io_out_bits_wstrb_5),
    .io_out_bits_wstrb_6(wdataMux_io_out_bits_wstrb_6),
    .io_out_bits_wstrb_7(wdataMux_io_out_bits_wstrb_7),
    .io_out_bits_wstrb_8(wdataMux_io_out_bits_wstrb_8),
    .io_out_bits_wstrb_9(wdataMux_io_out_bits_wstrb_9),
    .io_out_bits_wstrb_10(wdataMux_io_out_bits_wstrb_10),
    .io_out_bits_wstrb_11(wdataMux_io_out_bits_wstrb_11),
    .io_out_bits_wstrb_12(wdataMux_io_out_bits_wstrb_12),
    .io_out_bits_wstrb_13(wdataMux_io_out_bits_wstrb_13),
    .io_out_bits_wstrb_14(wdataMux_io_out_bits_wstrb_14),
    .io_out_bits_wstrb_15(wdataMux_io_out_bits_wstrb_15),
    .io_out_bits_wstrb_16(wdataMux_io_out_bits_wstrb_16),
    .io_out_bits_wstrb_17(wdataMux_io_out_bits_wstrb_17),
    .io_out_bits_wstrb_18(wdataMux_io_out_bits_wstrb_18),
    .io_out_bits_wstrb_19(wdataMux_io_out_bits_wstrb_19),
    .io_out_bits_wstrb_20(wdataMux_io_out_bits_wstrb_20),
    .io_out_bits_wstrb_21(wdataMux_io_out_bits_wstrb_21),
    .io_out_bits_wstrb_22(wdataMux_io_out_bits_wstrb_22),
    .io_out_bits_wstrb_23(wdataMux_io_out_bits_wstrb_23),
    .io_out_bits_wstrb_24(wdataMux_io_out_bits_wstrb_24),
    .io_out_bits_wstrb_25(wdataMux_io_out_bits_wstrb_25),
    .io_out_bits_wstrb_26(wdataMux_io_out_bits_wstrb_26),
    .io_out_bits_wstrb_27(wdataMux_io_out_bits_wstrb_27),
    .io_out_bits_wstrb_28(wdataMux_io_out_bits_wstrb_28),
    .io_out_bits_wstrb_29(wdataMux_io_out_bits_wstrb_29),
    .io_out_bits_wstrb_30(wdataMux_io_out_bits_wstrb_30),
    .io_out_bits_wstrb_31(wdataMux_io_out_bits_wstrb_31),
    .io_out_bits_wstrb_32(wdataMux_io_out_bits_wstrb_32),
    .io_out_bits_wstrb_33(wdataMux_io_out_bits_wstrb_33),
    .io_out_bits_wstrb_34(wdataMux_io_out_bits_wstrb_34),
    .io_out_bits_wstrb_35(wdataMux_io_out_bits_wstrb_35),
    .io_out_bits_wstrb_36(wdataMux_io_out_bits_wstrb_36),
    .io_out_bits_wstrb_37(wdataMux_io_out_bits_wstrb_37),
    .io_out_bits_wstrb_38(wdataMux_io_out_bits_wstrb_38),
    .io_out_bits_wstrb_39(wdataMux_io_out_bits_wstrb_39),
    .io_out_bits_wstrb_40(wdataMux_io_out_bits_wstrb_40),
    .io_out_bits_wstrb_41(wdataMux_io_out_bits_wstrb_41),
    .io_out_bits_wstrb_42(wdataMux_io_out_bits_wstrb_42),
    .io_out_bits_wstrb_43(wdataMux_io_out_bits_wstrb_43),
    .io_out_bits_wstrb_44(wdataMux_io_out_bits_wstrb_44),
    .io_out_bits_wstrb_45(wdataMux_io_out_bits_wstrb_45),
    .io_out_bits_wstrb_46(wdataMux_io_out_bits_wstrb_46),
    .io_out_bits_wstrb_47(wdataMux_io_out_bits_wstrb_47),
    .io_out_bits_wstrb_48(wdataMux_io_out_bits_wstrb_48),
    .io_out_bits_wstrb_49(wdataMux_io_out_bits_wstrb_49),
    .io_out_bits_wstrb_50(wdataMux_io_out_bits_wstrb_50),
    .io_out_bits_wstrb_51(wdataMux_io_out_bits_wstrb_51),
    .io_out_bits_wstrb_52(wdataMux_io_out_bits_wstrb_52),
    .io_out_bits_wstrb_53(wdataMux_io_out_bits_wstrb_53),
    .io_out_bits_wstrb_54(wdataMux_io_out_bits_wstrb_54),
    .io_out_bits_wstrb_55(wdataMux_io_out_bits_wstrb_55),
    .io_out_bits_wstrb_56(wdataMux_io_out_bits_wstrb_56),
    .io_out_bits_wstrb_57(wdataMux_io_out_bits_wstrb_57),
    .io_out_bits_wstrb_58(wdataMux_io_out_bits_wstrb_58),
    .io_out_bits_wstrb_59(wdataMux_io_out_bits_wstrb_59),
    .io_out_bits_wstrb_60(wdataMux_io_out_bits_wstrb_60),
    .io_out_bits_wstrb_61(wdataMux_io_out_bits_wstrb_61),
    .io_out_bits_wstrb_62(wdataMux_io_out_bits_wstrb_62),
    .io_out_bits_wstrb_63(wdataMux_io_out_bits_wstrb_63)
  );
  MuxN_4 cmdDeqValidMux (
    .io_ins_0(cmdDeqValidMux_io_ins_0),
    .io_ins_1(cmdDeqValidMux_io_ins_1),
    .io_sel(cmdDeqValidMux_io_sel),
    .io_out(cmdDeqValidMux_io_out)
  );
  MuxN_8 dramCmdMux (
    .io_ins_0_valid(dramCmdMux_io_ins_0_valid),
    .io_ins_0_bits_addr(dramCmdMux_io_ins_0_bits_addr),
    .io_ins_0_bits_size(dramCmdMux_io_ins_0_bits_size),
    .io_ins_0_bits_isWr(dramCmdMux_io_ins_0_bits_isWr),
    .io_ins_0_bits_tag_uid(dramCmdMux_io_ins_0_bits_tag_uid),
    .io_ins_0_bits_tag_streamId(dramCmdMux_io_ins_0_bits_tag_streamId),
    .io_ins_1_valid(dramCmdMux_io_ins_1_valid),
    .io_ins_1_bits_addr(dramCmdMux_io_ins_1_bits_addr),
    .io_ins_1_bits_size(dramCmdMux_io_ins_1_bits_size),
    .io_ins_1_bits_isWr(dramCmdMux_io_ins_1_bits_isWr),
    .io_ins_1_bits_tag_uid(dramCmdMux_io_ins_1_bits_tag_uid),
    .io_ins_1_bits_tag_streamId(dramCmdMux_io_ins_1_bits_tag_streamId),
    .io_sel(dramCmdMux_io_sel),
    .io_out_valid(dramCmdMux_io_out_valid),
    .io_out_bits_addr(dramCmdMux_io_out_bits_addr),
    .io_out_bits_size(dramCmdMux_io_out_bits_size),
    .io_out_bits_isWr(dramCmdMux_io_out_bits_isWr),
    .io_out_bits_tag_uid(dramCmdMux_io_out_bits_tag_uid),
    .io_out_bits_tag_streamId(dramCmdMux_io_out_bits_tag_streamId)
  );
  FF_143 FF_1 (
    .clock(FF_1_clock),
    .reset(FF_1_reset),
    .io_in(FF_1_io_in),
    .io_out(FF_1_io_out),
    .io_enable(FF_1_io_enable)
  );
  FF_136 FF_2 (
    .clock(FF_2_clock),
    .reset(FF_2_reset),
    .io_in(FF_2_io_in),
    .io_init(FF_2_io_init),
    .io_reset(FF_2_io_reset),
    .io_out(FF_2_io_out),
    .io_enable(FF_2_io_enable)
  );
  FF_145 FF_3 (
    .clock(FF_3_clock),
    .reset(FF_3_reset),
    .io_in(FF_3_io_in),
    .io_out(FF_3_io_out),
    .io_enable(FF_3_io_enable)
  );
  FF_115 FF_4 (
    .clock(FF_4_clock),
    .reset(FF_4_reset),
    .io_in(FF_4_io_in),
    .io_init(FF_4_io_init),
    .io_reset(FF_4_io_reset),
    .io_out(FF_4_io_out),
    .io_enable(FF_4_io_enable)
  );
  FF_137 FF_5 (
    .clock(FF_5_clock),
    .reset(FF_5_reset),
    .io_in(FF_5_io_in),
    .io_out(FF_5_io_out),
    .io_enable(FF_5_io_enable)
  );
  MuxN_5 wrespReadyMux (
    .io_ins_0(wrespReadyMux_io_ins_0),
    .io_out(wrespReadyMux_io_out)
  );
  MuxN_4 gatherLoadIssueMux (
    .io_ins_0(gatherLoadIssueMux_io_ins_0),
    .io_ins_1(gatherLoadIssueMux_io_ins_1),
    .io_sel(gatherLoadIssueMux_io_sel),
    .io_out(gatherLoadIssueMux_io_out)
  );
  Counter_18 gatherLoadIssue (
    .clock(gatherLoadIssue_clock),
    .reset(gatherLoadIssue_reset),
    .io_out(gatherLoadIssue_io_out),
    .io_reset(gatherLoadIssue_io_reset),
    .io_enable(gatherLoadIssue_io_enable)
  );
  MuxN_4 gatherLoadSkipMux (
    .io_ins_0(gatherLoadSkipMux_io_ins_0),
    .io_ins_1(gatherLoadSkipMux_io_ins_1),
    .io_sel(gatherLoadSkipMux_io_sel),
    .io_out(gatherLoadSkipMux_io_out)
  );
  Counter_18 gatherLoadSkip (
    .clock(gatherLoadSkip_clock),
    .reset(gatherLoadSkip_reset),
    .io_out(gatherLoadSkip_io_out),
    .io_reset(gatherLoadSkip_io_reset),
    .io_enable(gatherLoadSkip_io_enable)
  );
  MuxN_4 scatterLoadIssueMux (
    .io_ins_0(scatterLoadIssueMux_io_ins_0),
    .io_ins_1(scatterLoadIssueMux_io_ins_1),
    .io_sel(scatterLoadIssueMux_io_sel),
    .io_out(scatterLoadIssueMux_io_out)
  );
  Counter_18 scatterLoadIssue (
    .clock(scatterLoadIssue_clock),
    .reset(scatterLoadIssue_reset),
    .io_out(scatterLoadIssue_io_out),
    .io_reset(scatterLoadIssue_io_reset),
    .io_enable(scatterLoadIssue_io_enable)
  );
  MuxN_4 scatterLoadSkipMux (
    .io_ins_0(scatterLoadSkipMux_io_ins_0),
    .io_ins_1(scatterLoadSkipMux_io_ins_1),
    .io_sel(scatterLoadSkipMux_io_sel),
    .io_out(scatterLoadSkipMux_io_out)
  );
  Counter_18 scatterLoadSkip (
    .clock(scatterLoadSkip_clock),
    .reset(scatterLoadSkip_reset),
    .io_out(scatterLoadSkip_io_out),
    .io_reset(scatterLoadSkip_io_reset),
    .io_enable(scatterLoadSkip_io_enable)
  );
  MuxN_4 scatterStoreIssueMux (
    .io_ins_0(scatterStoreIssueMux_io_ins_0),
    .io_ins_1(scatterStoreIssueMux_io_ins_1),
    .io_sel(scatterStoreIssueMux_io_sel),
    .io_out(scatterStoreIssueMux_io_out)
  );
  Counter_18 scatterStoreIssue (
    .clock(scatterStoreIssue_clock),
    .reset(scatterStoreIssue_reset),
    .io_out(scatterStoreIssue_io_out),
    .io_reset(scatterStoreIssue_io_reset),
    .io_enable(scatterStoreIssue_io_enable)
  );
  MuxN_4 scatterStoreSkipMux (
    .io_ins_0(scatterStoreSkipMux_io_ins_0),
    .io_ins_1(scatterStoreSkipMux_io_ins_1),
    .io_sel(scatterStoreSkipMux_io_sel),
    .io_out(scatterStoreSkipMux_io_out)
  );
  Counter_18 scatterStoreSkip (
    .clock(scatterStoreSkip_clock),
    .reset(scatterStoreSkip_reset),
    .io_out(scatterStoreSkip_io_out),
    .io_reset(scatterStoreSkip_io_reset),
    .io_enable(scatterStoreSkip_io_enable)
  );
  FIFOWidthConvert denseLoadBuffers_0 (
    .clock(denseLoadBuffers_0_clock),
    .reset(denseLoadBuffers_0_reset),
    .io_enq_0(denseLoadBuffers_0_io_enq_0),
    .io_enq_1(denseLoadBuffers_0_io_enq_1),
    .io_enq_2(denseLoadBuffers_0_io_enq_2),
    .io_enq_3(denseLoadBuffers_0_io_enq_3),
    .io_enq_4(denseLoadBuffers_0_io_enq_4),
    .io_enq_5(denseLoadBuffers_0_io_enq_5),
    .io_enq_6(denseLoadBuffers_0_io_enq_6),
    .io_enq_7(denseLoadBuffers_0_io_enq_7),
    .io_enq_8(denseLoadBuffers_0_io_enq_8),
    .io_enq_9(denseLoadBuffers_0_io_enq_9),
    .io_enq_10(denseLoadBuffers_0_io_enq_10),
    .io_enq_11(denseLoadBuffers_0_io_enq_11),
    .io_enq_12(denseLoadBuffers_0_io_enq_12),
    .io_enq_13(denseLoadBuffers_0_io_enq_13),
    .io_enq_14(denseLoadBuffers_0_io_enq_14),
    .io_enq_15(denseLoadBuffers_0_io_enq_15),
    .io_enqVld(denseLoadBuffers_0_io_enqVld),
    .io_deq_0(denseLoadBuffers_0_io_deq_0),
    .io_deqVld(denseLoadBuffers_0_io_deqVld),
    .io_full(denseLoadBuffers_0_io_full),
    .io_empty(denseLoadBuffers_0_io_empty),
    .io_almostEmpty(denseLoadBuffers_0_io_almostEmpty),
    .io_almostFull(denseLoadBuffers_0_io_almostFull)
  );
  Counter_18 Counter (
    .clock(Counter_clock),
    .reset(Counter_reset),
    .io_out(Counter_io_out),
    .io_reset(Counter_io_reset),
    .io_enable(Counter_io_enable)
  );
  Counter_18 Counter_1 (
    .clock(Counter_1_clock),
    .reset(Counter_1_reset),
    .io_out(Counter_1_io_out),
    .io_reset(Counter_1_io_reset),
    .io_enable(Counter_1_io_enable)
  );
  Counter_18 Counter_2 (
    .clock(Counter_2_clock),
    .reset(Counter_2_reset),
    .io_out(Counter_2_io_out),
    .io_reset(Counter_2_io_reset),
    .io_enable(Counter_2_io_enable)
  );
  Counter_18 Counter_3 (
    .clock(Counter_3_clock),
    .reset(Counter_3_reset),
    .io_out(Counter_3_io_out),
    .io_reset(Counter_3_io_reset),
    .io_enable(Counter_3_io_enable)
  );
  Counter_18 Counter_4 (
    .clock(Counter_4_clock),
    .reset(Counter_4_reset),
    .io_out(Counter_4_io_out),
    .io_reset(Counter_4_io_reset),
    .io_enable(Counter_4_io_enable)
  );
  SRFF SRFF (
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output_data(SRFF_io_output_data)
  );
  SRFF SRFF_1 (
    .clock(SRFF_1_clock),
    .reset(SRFF_1_reset),
    .io_input_set(SRFF_1_io_input_set),
    .io_input_reset(SRFF_1_io_input_reset),
    .io_input_asyn_reset(SRFF_1_io_input_asyn_reset),
    .io_output_data(SRFF_1_io_output_data)
  );
  FF_145 FF_6 (
    .clock(FF_6_clock),
    .reset(FF_6_reset),
    .io_in(FF_6_io_in),
    .io_out(FF_6_io_out),
    .io_enable(FF_6_io_enable)
  );
  FF_180 FF_7 (
    .clock(FF_7_clock),
    .reset(FF_7_reset),
    .io_in(FF_7_io_in),
    .io_out(FF_7_io_out),
    .io_enable(FF_7_io_enable)
  );
  FIFOWidthConvert_1 denseStoreBuffers_0 (
    .clock(denseStoreBuffers_0_clock),
    .reset(denseStoreBuffers_0_reset),
    .io_enqVld(denseStoreBuffers_0_io_enqVld),
    .io_deq_0(denseStoreBuffers_0_io_deq_0),
    .io_deq_1(denseStoreBuffers_0_io_deq_1),
    .io_deq_2(denseStoreBuffers_0_io_deq_2),
    .io_deq_3(denseStoreBuffers_0_io_deq_3),
    .io_deq_4(denseStoreBuffers_0_io_deq_4),
    .io_deq_5(denseStoreBuffers_0_io_deq_5),
    .io_deq_6(denseStoreBuffers_0_io_deq_6),
    .io_deq_7(denseStoreBuffers_0_io_deq_7),
    .io_deq_8(denseStoreBuffers_0_io_deq_8),
    .io_deq_9(denseStoreBuffers_0_io_deq_9),
    .io_deq_10(denseStoreBuffers_0_io_deq_10),
    .io_deq_11(denseStoreBuffers_0_io_deq_11),
    .io_deq_12(denseStoreBuffers_0_io_deq_12),
    .io_deq_13(denseStoreBuffers_0_io_deq_13),
    .io_deq_14(denseStoreBuffers_0_io_deq_14),
    .io_deq_15(denseStoreBuffers_0_io_deq_15),
    .io_deqStrb(denseStoreBuffers_0_io_deqStrb),
    .io_deqVld(denseStoreBuffers_0_io_deqVld),
    .io_full(denseStoreBuffers_0_io_full),
    .io_empty(denseStoreBuffers_0_io_empty),
    .io_almostEmpty(denseStoreBuffers_0_io_almostEmpty),
    .io_almostFull(denseStoreBuffers_0_io_almostFull)
  );
  Counter_15 Counter_5 (
    .clock(Counter_5_clock),
    .reset(Counter_5_reset),
    .io_max(Counter_5_io_max),
    .io_stride(Counter_5_io_stride),
    .io_out(Counter_5_io_out),
    .io_last(Counter_5_io_last),
    .io_reset(Counter_5_io_reset),
    .io_enable(Counter_5_io_enable),
    .io_done(Counter_5_io_done)
  );
  FF_137 FF_8 (
    .clock(FF_8_clock),
    .reset(FF_8_reset),
    .io_in(FF_8_io_in),
    .io_out(FF_8_io_out),
    .io_enable(FF_8_io_enable)
  );
  FIFOCounter FIFOCounter (
    .clock(FIFOCounter_clock),
    .reset(FIFOCounter_reset),
    .io_enqVld(FIFOCounter_io_enqVld),
    .io_full(FIFOCounter_io_full),
    .io_empty(FIFOCounter_io_empty)
  );
  Counter_18 Counter_6 (
    .clock(Counter_6_clock),
    .reset(Counter_6_reset),
    .io_out(Counter_6_io_out),
    .io_reset(Counter_6_io_reset),
    .io_enable(Counter_6_io_enable)
  );
  Counter_18 Counter_7 (
    .clock(Counter_7_clock),
    .reset(Counter_7_reset),
    .io_out(Counter_7_io_out),
    .io_reset(Counter_7_io_reset),
    .io_enable(Counter_7_io_enable)
  );
  Counter_18 Counter_8 (
    .clock(Counter_8_clock),
    .reset(Counter_8_reset),
    .io_out(Counter_8_io_out),
    .io_reset(Counter_8_io_reset),
    .io_enable(Counter_8_io_enable)
  );
  FF_145 burstCounterMaxLatch (
    .clock(burstCounterMaxLatch_clock),
    .reset(burstCounterMaxLatch_reset),
    .io_in(burstCounterMaxLatch_io_in),
    .io_out(burstCounterMaxLatch_io_out),
    .io_enable(burstCounterMaxLatch_io_enable)
  );
  FF_115 dramReadyFF (
    .clock(dramReadyFF_clock),
    .reset(dramReadyFF_reset),
    .io_in(dramReadyFF_io_in),
    .io_init(dramReadyFF_io_init),
    .io_reset(dramReadyFF_io_reset),
    .io_out(dramReadyFF_io_out),
    .io_enable(dramReadyFF_io_enable)
  );
  Counter_18 cycleCount (
    .clock(cycleCount_clock),
    .reset(cycleCount_reset),
    .io_out(cycleCount_io_out),
    .io_reset(cycleCount_io_reset),
    .io_enable(cycleCount_io_enable)
  );
  Counter_18 rdataEnqCount (
    .clock(rdataEnqCount_clock),
    .reset(rdataEnqCount_reset),
    .io_out(rdataEnqCount_io_out),
    .io_reset(rdataEnqCount_io_reset),
    .io_enable(rdataEnqCount_io_enable)
  );
  Counter_18 wdataCount (
    .clock(wdataCount_clock),
    .reset(wdataCount_reset),
    .io_out(wdataCount_io_out),
    .io_reset(wdataCount_io_reset),
    .io_enable(wdataCount_io_enable)
  );
  Counter_18 Counter_9 (
    .clock(Counter_9_clock),
    .reset(Counter_9_reset),
    .io_out(Counter_9_io_out),
    .io_reset(Counter_9_io_reset),
    .io_enable(Counter_9_io_enable)
  );
  Counter_18 Counter_10 (
    .clock(Counter_10_clock),
    .reset(Counter_10_reset),
    .io_out(Counter_10_io_out),
    .io_reset(Counter_10_io_reset),
    .io_enable(Counter_10_io_enable)
  );
  Counter_18 Counter_11 (
    .clock(Counter_11_clock),
    .reset(Counter_11_reset),
    .io_out(Counter_11_io_out),
    .io_reset(Counter_11_io_reset),
    .io_enable(Counter_11_io_enable)
  );
  Counter_18 Counter_12 (
    .clock(Counter_12_clock),
    .reset(Counter_12_reset),
    .io_out(Counter_12_io_out),
    .io_reset(Counter_12_io_reset),
    .io_enable(Counter_12_io_enable)
  );
  Counter_18 Counter_13 (
    .clock(Counter_13_clock),
    .reset(Counter_13_reset),
    .io_out(Counter_13_io_out),
    .io_reset(Counter_13_io_reset),
    .io_enable(Counter_13_io_enable)
  );
  Counter_18 Counter_14 (
    .clock(Counter_14_clock),
    .reset(Counter_14_reset),
    .io_out(Counter_14_io_out),
    .io_reset(Counter_14_io_reset),
    .io_enable(Counter_14_io_enable)
  );
  Counter_18 Counter_15 (
    .clock(Counter_15_clock),
    .reset(Counter_15_reset),
    .io_out(Counter_15_io_out),
    .io_reset(Counter_15_io_reset),
    .io_enable(Counter_15_io_enable)
  );
  Counter_18 Counter_16 (
    .clock(Counter_16_clock),
    .reset(Counter_16_reset),
    .io_out(Counter_16_io_out),
    .io_reset(Counter_16_io_reset),
    .io_enable(Counter_16_io_enable)
  );
  Counter_18 Counter_17 (
    .clock(Counter_17_clock),
    .reset(Counter_17_reset),
    .io_out(Counter_17_io_out),
    .io_reset(Counter_17_io_reset),
    .io_enable(Counter_17_io_enable)
  );
  Counter_18 Counter_18 (
    .clock(Counter_18_clock),
    .reset(Counter_18_reset),
    .io_out(Counter_18_io_out),
    .io_reset(Counter_18_io_reset),
    .io_enable(Counter_18_io_enable)
  );
  Counter_18 Counter_19 (
    .clock(Counter_19_clock),
    .reset(Counter_19_reset),
    .io_out(Counter_19_io_out),
    .io_reset(Counter_19_io_reset),
    .io_enable(Counter_19_io_enable)
  );
  Counter_18 Counter_20 (
    .clock(Counter_20_clock),
    .reset(Counter_20_reset),
    .io_out(Counter_20_io_out),
    .io_reset(Counter_20_io_reset),
    .io_enable(Counter_20_io_enable)
  );
  Counter_18 Counter_21 (
    .clock(Counter_21_clock),
    .reset(Counter_21_reset),
    .io_out(Counter_21_io_out),
    .io_reset(Counter_21_io_reset),
    .io_enable(Counter_21_io_enable)
  );
  Counter_18 Counter_22 (
    .clock(Counter_22_clock),
    .reset(Counter_22_reset),
    .io_out(Counter_22_io_out),
    .io_reset(Counter_22_io_reset),
    .io_enable(Counter_22_io_enable)
  );
  Counter_18 Counter_23 (
    .clock(Counter_23_clock),
    .reset(Counter_23_reset),
    .io_out(Counter_23_io_out),
    .io_reset(Counter_23_io_reset),
    .io_enable(Counter_23_io_enable)
  );
  Counter_18 Counter_24 (
    .clock(Counter_24_clock),
    .reset(Counter_24_reset),
    .io_out(Counter_24_io_out),
    .io_reset(Counter_24_io_reset),
    .io_enable(Counter_24_io_enable)
  );
  Counter_18 Counter_25 (
    .clock(Counter_25_clock),
    .reset(Counter_25_reset),
    .io_out(Counter_25_io_out),
    .io_reset(Counter_25_io_reset),
    .io_enable(Counter_25_io_enable)
  );
  Counter_18 Counter_26 (
    .clock(Counter_26_clock),
    .reset(Counter_26_reset),
    .io_out(Counter_26_io_out),
    .io_reset(Counter_26_io_reset),
    .io_enable(Counter_26_io_enable)
  );
  Counter_18 Counter_27 (
    .clock(Counter_27_clock),
    .reset(Counter_27_reset),
    .io_out(Counter_27_io_out),
    .io_reset(Counter_27_io_reset),
    .io_enable(Counter_27_io_enable)
  );
  Counter_18 Counter_28 (
    .clock(Counter_28_clock),
    .reset(Counter_28_reset),
    .io_out(Counter_28_io_out),
    .io_reset(Counter_28_io_reset),
    .io_enable(Counter_28_io_enable)
  );
  Counter_18 Counter_29 (
    .clock(Counter_29_clock),
    .reset(Counter_29_reset),
    .io_out(Counter_29_io_out),
    .io_reset(Counter_29_io_reset),
    .io_enable(Counter_29_io_enable)
  );
  Counter_18 Counter_30 (
    .clock(Counter_30_clock),
    .reset(Counter_30_reset),
    .io_out(Counter_30_io_out),
    .io_reset(Counter_30_io_reset),
    .io_enable(Counter_30_io_enable)
  );
  Counter_18 Counter_31 (
    .clock(Counter_31_clock),
    .reset(Counter_31_reset),
    .io_out(Counter_31_io_out),
    .io_reset(Counter_31_io_reset),
    .io_enable(Counter_31_io_enable)
  );
  Counter_18 Counter_32 (
    .clock(Counter_32_clock),
    .reset(Counter_32_reset),
    .io_out(Counter_32_io_out),
    .io_reset(Counter_32_io_reset),
    .io_enable(Counter_32_io_enable)
  );
  Counter_18 Counter_33 (
    .clock(Counter_33_clock),
    .reset(Counter_33_reset),
    .io_out(Counter_33_io_out),
    .io_reset(Counter_33_io_reset),
    .io_enable(Counter_33_io_enable)
  );
  Counter_18 Counter_34 (
    .clock(Counter_34_clock),
    .reset(Counter_34_reset),
    .io_out(Counter_34_io_out),
    .io_reset(Counter_34_io_reset),
    .io_enable(Counter_34_io_enable)
  );
  FF_143 FF_9 (
    .clock(FF_9_clock),
    .reset(FF_9_reset),
    .io_in(FF_9_io_in),
    .io_out(FF_9_io_out),
    .io_enable(FF_9_io_enable)
  );
  Counter_18 Counter_35 (
    .clock(Counter_35_clock),
    .reset(Counter_35_reset),
    .io_out(Counter_35_io_out),
    .io_reset(Counter_35_io_reset),
    .io_enable(Counter_35_io_enable)
  );
  Counter_18 Counter_36 (
    .clock(Counter_36_clock),
    .reset(Counter_36_reset),
    .io_out(Counter_36_io_out),
    .io_reset(Counter_36_io_reset),
    .io_enable(Counter_36_io_enable)
  );
  Counter_18 Counter_37 (
    .clock(Counter_37_clock),
    .reset(Counter_37_reset),
    .io_out(Counter_37_io_out),
    .io_reset(Counter_37_io_reset),
    .io_enable(Counter_37_io_enable)
  );
  Counter_18 Counter_38 (
    .clock(Counter_38_clock),
    .reset(Counter_38_reset),
    .io_out(Counter_38_io_out),
    .io_reset(Counter_38_io_reset),
    .io_enable(Counter_38_io_enable)
  );
  Counter_18 Counter_39 (
    .clock(Counter_39_clock),
    .reset(Counter_39_reset),
    .io_out(Counter_39_io_out),
    .io_reset(Counter_39_io_reset),
    .io_enable(Counter_39_io_enable)
  );
  Counter_18 Counter_40 (
    .clock(Counter_40_clock),
    .reset(Counter_40_reset),
    .io_out(Counter_40_io_out),
    .io_reset(Counter_40_io_reset),
    .io_enable(Counter_40_io_enable)
  );
  Counter_18 Counter_41 (
    .clock(Counter_41_clock),
    .reset(Counter_41_reset),
    .io_out(Counter_41_io_out),
    .io_reset(Counter_41_io_reset),
    .io_enable(Counter_41_io_enable)
  );
  Counter_18 Counter_42 (
    .clock(Counter_42_clock),
    .reset(Counter_42_reset),
    .io_out(Counter_42_io_out),
    .io_reset(Counter_42_io_reset),
    .io_enable(Counter_42_io_enable)
  );
  Counter_18 Counter_43 (
    .clock(Counter_43_clock),
    .reset(Counter_43_reset),
    .io_out(Counter_43_io_out),
    .io_reset(Counter_43_io_reset),
    .io_enable(Counter_43_io_enable)
  );
  Counter_18 Counter_44 (
    .clock(Counter_44_clock),
    .reset(Counter_44_reset),
    .io_out(Counter_44_io_out),
    .io_reset(Counter_44_io_reset),
    .io_enable(Counter_44_io_enable)
  );
  Counter_18 Counter_45 (
    .clock(Counter_45_clock),
    .reset(Counter_45_reset),
    .io_out(Counter_45_io_out),
    .io_reset(Counter_45_io_reset),
    .io_enable(Counter_45_io_enable)
  );
  Counter_18 Counter_46 (
    .clock(Counter_46_clock),
    .reset(Counter_46_reset),
    .io_out(Counter_46_io_out),
    .io_reset(Counter_46_io_reset),
    .io_enable(Counter_46_io_enable)
  );
  Counter_18 Counter_47 (
    .clock(Counter_47_clock),
    .reset(Counter_47_reset),
    .io_out(Counter_47_io_out),
    .io_reset(Counter_47_io_reset),
    .io_enable(Counter_47_io_enable)
  );
  Counter_18 Counter_48 (
    .clock(Counter_48_clock),
    .reset(Counter_48_reset),
    .io_out(Counter_48_io_out),
    .io_reset(Counter_48_io_reset),
    .io_enable(Counter_48_io_enable)
  );
  Counter_18 Counter_49 (
    .clock(Counter_49_clock),
    .reset(Counter_49_reset),
    .io_out(Counter_49_io_out),
    .io_reset(Counter_49_io_reset),
    .io_enable(Counter_49_io_enable)
  );
  Counter_18 Counter_50 (
    .clock(Counter_50_clock),
    .reset(Counter_50_reset),
    .io_out(Counter_50_io_out),
    .io_reset(Counter_50_io_reset),
    .io_enable(Counter_50_io_enable)
  );
  Counter_18 Counter_51 (
    .clock(Counter_51_clock),
    .reset(Counter_51_reset),
    .io_out(Counter_51_io_out),
    .io_reset(Counter_51_io_reset),
    .io_enable(Counter_51_io_enable)
  );
  Counter_18 Counter_52 (
    .clock(Counter_52_clock),
    .reset(Counter_52_reset),
    .io_out(Counter_52_io_out),
    .io_reset(Counter_52_io_reset),
    .io_enable(Counter_52_io_enable)
  );
  Counter_18 Counter_53 (
    .clock(Counter_53_clock),
    .reset(Counter_53_reset),
    .io_out(Counter_53_io_out),
    .io_reset(Counter_53_io_reset),
    .io_enable(Counter_53_io_enable)
  );
  Counter_18 Counter_54 (
    .clock(Counter_54_clock),
    .reset(Counter_54_reset),
    .io_out(Counter_54_io_out),
    .io_reset(Counter_54_io_reset),
    .io_enable(Counter_54_io_enable)
  );
  Counter_18 Counter_55 (
    .clock(Counter_55_clock),
    .reset(Counter_55_reset),
    .io_out(Counter_55_io_out),
    .io_reset(Counter_55_io_reset),
    .io_enable(Counter_55_io_enable)
  );
  Counter_18 Counter_56 (
    .clock(Counter_56_clock),
    .reset(Counter_56_reset),
    .io_out(Counter_56_io_out),
    .io_reset(Counter_56_io_reset),
    .io_enable(Counter_56_io_enable)
  );
  Counter_18 Counter_57 (
    .clock(Counter_57_clock),
    .reset(Counter_57_reset),
    .io_out(Counter_57_io_out),
    .io_reset(Counter_57_io_reset),
    .io_enable(Counter_57_io_enable)
  );
  Counter_18 Counter_58 (
    .clock(Counter_58_clock),
    .reset(Counter_58_reset),
    .io_out(Counter_58_io_out),
    .io_reset(Counter_58_io_reset),
    .io_enable(Counter_58_io_enable)
  );
  Counter_18 Counter_59 (
    .clock(Counter_59_clock),
    .reset(Counter_59_reset),
    .io_out(Counter_59_io_out),
    .io_reset(Counter_59_io_reset),
    .io_enable(Counter_59_io_enable)
  );
  FF_136 FF_10 (
    .clock(FF_10_clock),
    .reset(FF_10_reset),
    .io_in(FF_10_io_in),
    .io_init(FF_10_io_init),
    .io_reset(FF_10_io_reset),
    .io_out(FF_10_io_out),
    .io_enable(FF_10_io_enable)
  );
  FF_265 FF_11 (
    .clock(FF_11_clock),
    .reset(FF_11_reset),
    .io_in(FF_11_io_in),
    .io_out(FF_11_io_out),
    .io_enable(FF_11_io_enable)
  );
  FF_266 FF_12 (
    .clock(FF_12_clock),
    .reset(FF_12_reset),
    .io_in(FF_12_io_in),
    .io_out(FF_12_io_out),
    .io_enable(FF_12_io_enable)
  );
  FF_115 FF_13 (
    .clock(FF_13_clock),
    .reset(FF_13_reset),
    .io_in(FF_13_io_in),
    .io_init(FF_13_io_init),
    .io_reset(FF_13_io_reset),
    .io_out(FF_13_io_out),
    .io_enable(FF_13_io_enable)
  );
  FF_268 FF_14 (
    .clock(FF_14_clock),
    .reset(FF_14_reset),
    .io_in(FF_14_io_in),
    .io_out(FF_14_io_out),
    .io_enable(FF_14_io_enable)
  );
  FF_136 FF_15 (
    .clock(FF_15_clock),
    .reset(FF_15_reset),
    .io_in(FF_15_io_in),
    .io_init(FF_15_io_init),
    .io_reset(FF_15_io_reset),
    .io_out(FF_15_io_out),
    .io_enable(FF_15_io_enable)
  );
  FF_265 FF_16 (
    .clock(FF_16_clock),
    .reset(FF_16_reset),
    .io_in(FF_16_io_in),
    .io_out(FF_16_io_out),
    .io_enable(FF_16_io_enable)
  );
  FF_180 FF_17 (
    .clock(FF_17_clock),
    .reset(FF_17_reset),
    .io_in(FF_17_io_in),
    .io_out(FF_17_io_out),
    .io_enable(FF_17_io_enable)
  );
  FF_136 FF_18 (
    .clock(FF_18_clock),
    .reset(FF_18_reset),
    .io_in(FF_18_io_in),
    .io_init(FF_18_io_init),
    .io_reset(FF_18_io_reset),
    .io_out(FF_18_io_out),
    .io_enable(FF_18_io_enable)
  );
  FF_180 FF_19 (
    .clock(FF_19_clock),
    .reset(FF_19_reset),
    .io_in(FF_19_io_in),
    .io_out(FF_19_io_out),
    .io_enable(FF_19_io_enable)
  );
  FF_136 FF_20 (
    .clock(FF_20_clock),
    .reset(FF_20_reset),
    .io_in(FF_20_io_in),
    .io_init(FF_20_io_init),
    .io_reset(FF_20_io_reset),
    .io_out(FF_20_io_out),
    .io_enable(FF_20_io_enable)
  );
  FF_180 FF_21 (
    .clock(FF_21_clock),
    .reset(FF_21_reset),
    .io_in(FF_21_io_in),
    .io_out(FF_21_io_out),
    .io_enable(FF_21_io_enable)
  );
  FF_136 FF_22 (
    .clock(FF_22_clock),
    .reset(FF_22_reset),
    .io_in(FF_22_io_in),
    .io_init(FF_22_io_init),
    .io_reset(FF_22_io_reset),
    .io_out(FF_22_io_out),
    .io_enable(FF_22_io_enable)
  );
  Counter_18 Counter_60 (
    .clock(Counter_60_clock),
    .reset(Counter_60_reset),
    .io_out(Counter_60_io_out),
    .io_reset(Counter_60_io_reset),
    .io_enable(Counter_60_io_enable)
  );
  Counter_18 Counter_61 (
    .clock(Counter_61_clock),
    .reset(Counter_61_reset),
    .io_out(Counter_61_io_out),
    .io_reset(Counter_61_io_reset),
    .io_enable(Counter_61_io_enable)
  );
  Counter_18 Counter_62 (
    .clock(Counter_62_clock),
    .reset(Counter_62_reset),
    .io_out(Counter_62_io_out),
    .io_reset(Counter_62_io_reset),
    .io_enable(Counter_62_io_enable)
  );
  Counter_18 Counter_63 (
    .clock(Counter_63_clock),
    .reset(Counter_63_reset),
    .io_out(Counter_63_io_out),
    .io_reset(Counter_63_io_reset),
    .io_enable(Counter_63_io_enable)
  );
  Counter_18 Counter_64 (
    .clock(Counter_64_clock),
    .reset(Counter_64_reset),
    .io_out(Counter_64_io_out),
    .io_reset(Counter_64_io_reset),
    .io_enable(Counter_64_io_enable)
  );
  Counter_18 Counter_65 (
    .clock(Counter_65_clock),
    .reset(Counter_65_reset),
    .io_out(Counter_65_io_out),
    .io_reset(Counter_65_io_reset),
    .io_enable(Counter_65_io_enable)
  );
  Counter_18 Counter_66 (
    .clock(Counter_66_clock),
    .reset(Counter_66_reset),
    .io_out(Counter_66_io_out),
    .io_reset(Counter_66_io_reset),
    .io_enable(Counter_66_io_enable)
  );
  Counter_18 Counter_67 (
    .clock(Counter_67_clock),
    .reset(Counter_67_reset),
    .io_out(Counter_67_io_out),
    .io_reset(Counter_67_io_reset),
    .io_enable(Counter_67_io_enable)
  );
  Counter_18 Counter_68 (
    .clock(Counter_68_clock),
    .reset(Counter_68_reset),
    .io_out(Counter_68_io_out),
    .io_reset(Counter_68_io_reset),
    .io_enable(Counter_68_io_enable)
  );
  Counter_18 Counter_69 (
    .clock(Counter_69_clock),
    .reset(Counter_69_reset),
    .io_out(Counter_69_io_out),
    .io_reset(Counter_69_io_reset),
    .io_enable(Counter_69_io_enable)
  );
  Counter_18 Counter_70 (
    .clock(Counter_70_clock),
    .reset(Counter_70_reset),
    .io_out(Counter_70_io_out),
    .io_reset(Counter_70_io_reset),
    .io_enable(Counter_70_io_enable)
  );
  Counter_18 Counter_71 (
    .clock(Counter_71_clock),
    .reset(Counter_71_reset),
    .io_out(Counter_71_io_out),
    .io_reset(Counter_71_io_reset),
    .io_enable(Counter_71_io_enable)
  );
  Counter_18 Counter_72 (
    .clock(Counter_72_clock),
    .reset(Counter_72_reset),
    .io_out(Counter_72_io_out),
    .io_reset(Counter_72_io_reset),
    .io_enable(Counter_72_io_enable)
  );
  FF_136 FF_23 (
    .clock(FF_23_clock),
    .reset(FF_23_reset),
    .io_in(FF_23_io_in),
    .io_init(FF_23_io_init),
    .io_reset(FF_23_io_reset),
    .io_out(FF_23_io_out),
    .io_enable(FF_23_io_enable)
  );
  FF_265 FF_24 (
    .clock(FF_24_clock),
    .reset(FF_24_reset),
    .io_in(FF_24_io_in),
    .io_out(FF_24_io_out),
    .io_enable(FF_24_io_enable)
  );
  FF_266 FF_25 (
    .clock(FF_25_clock),
    .reset(FF_25_reset),
    .io_in(FF_25_io_in),
    .io_out(FF_25_io_out),
    .io_enable(FF_25_io_enable)
  );
  FF_268 FF_26 (
    .clock(FF_26_clock),
    .reset(FF_26_reset),
    .io_in(FF_26_io_in),
    .io_out(FF_26_io_out),
    .io_enable(FF_26_io_enable)
  );
  FF_136 FF_27 (
    .clock(FF_27_clock),
    .reset(FF_27_reset),
    .io_in(FF_27_io_in),
    .io_init(FF_27_io_init),
    .io_reset(FF_27_io_reset),
    .io_out(FF_27_io_out),
    .io_enable(FF_27_io_enable)
  );
  FF_265 FF_28 (
    .clock(FF_28_clock),
    .reset(FF_28_reset),
    .io_in(FF_28_io_in),
    .io_out(FF_28_io_out),
    .io_enable(FF_28_io_enable)
  );
  FF_180 FF_29 (
    .clock(FF_29_clock),
    .reset(FF_29_reset),
    .io_in(FF_29_io_in),
    .io_out(FF_29_io_out),
    .io_enable(FF_29_io_enable)
  );
  FF_136 FF_30 (
    .clock(FF_30_clock),
    .reset(FF_30_reset),
    .io_in(FF_30_io_in),
    .io_init(FF_30_io_init),
    .io_reset(FF_30_io_reset),
    .io_out(FF_30_io_out),
    .io_enable(FF_30_io_enable)
  );
  FF_180 FF_31 (
    .clock(FF_31_clock),
    .reset(FF_31_reset),
    .io_in(FF_31_io_in),
    .io_out(FF_31_io_out),
    .io_enable(FF_31_io_enable)
  );
  FF_136 FF_32 (
    .clock(FF_32_clock),
    .reset(FF_32_reset),
    .io_in(FF_32_io_in),
    .io_init(FF_32_io_init),
    .io_reset(FF_32_io_reset),
    .io_out(FF_32_io_out),
    .io_enable(FF_32_io_enable)
  );
  FF_180 FF_33 (
    .clock(FF_33_clock),
    .reset(FF_33_reset),
    .io_in(FF_33_io_in),
    .io_out(FF_33_io_out),
    .io_enable(FF_33_io_enable)
  );
  FF_136 FF_34 (
    .clock(FF_34_clock),
    .reset(FF_34_reset),
    .io_in(FF_34_io_in),
    .io_init(FF_34_io_init),
    .io_reset(FF_34_io_reset),
    .io_out(FF_34_io_out),
    .io_enable(FF_34_io_enable)
  );
  assign _T_886 = io_app_loads_0_cmd_bits_addr[31:0];
  assign _T_887 = {32'h7f,_T_886};
  assign _T_891 = ~ cmdArbiter_io_full_0;
  assign _GEN_0 = {{48'd0}, sizeCounter_io_out};
  assign _T_894 = cmdArbiter_io_deq_0_addr + _GEN_0;
  assign _T_895 = _T_894[63:0];
  assign _T_896 = io_enable & cmdArbiter_io_deqReady;
  assign _T_897 = ~ cmdArbiter_io_deq_0_isWr;
  assign cmdRead = _T_896 & _T_897;
  assign cmdWrite = _T_896 & cmdArbiter_io_deq_0_isWr;
  assign _T_903 = isSparseMux_io_out ? 16'h1 : cmdArbiter_io_deq_0_size;
  assign _T_908 = isSparseMux_io_out ? 1'h0 : sizeCounter_io_done;
  assign _T_931 = cmdAddr_bits[63:6];
  assign _T_933 = {_T_931,6'h0};
  assign _T_938 = cmdArbiter_io_deq_0_size - sizeCounter_io_out;
  assign _T_939 = $unsigned(_T_938);
  assign _T_940 = _T_939[15:0];
  assign _T_942 = sizeCounter_io_done ? _T_940 : 16'h4000;
  assign _T_943 = isSparseMux_io_out ? cmdArbiter_io_deq_0_size : _T_942;
  assign _T_944 = _T_937_bits[15:6];
  assign _T_945 = _T_937_bits[5:0];
  assign _T_947 = _T_945 != 6'h0;
  assign _GEN_2 = {{9'd0}, _T_947};
  assign _T_948 = _T_944 + _GEN_2;
  assign _T_949 = _T_948[9:0];
  assign _T_950 = ~ dramCmdMux_io_out_bits_isWr;
  assign _T_951 = dramCmdMux_io_out_valid & _T_950;
  assign _T_978 = _T_971_bits[15:6];
  assign _T_979 = _T_971_bits[5:0];
  assign _T_981 = _T_979 != 6'h0;
  assign _GEN_3 = {{9'd0}, _T_981};
  assign _T_982 = _T_978 + _GEN_3;
  assign _T_983 = _T_982[9:0];
  assign _T_1027 = io_dram_rresp_bits_tag_streamId == 6'h0;
  assign _T_1028 = io_dram_rresp_valid & _T_1027;
  assign _T_1029 = ~ denseLoadBuffers_0_io_full;
  assign _T_1031 = ~ denseLoadBuffers_0_io_empty;
  assign _T_1046 = _T_1031 & io_app_loads_0_rdata_ready;
  assign _T_1051 = denseLoadBuffers_0_io_empty & denseLoadBuffers_0_io_deqVld;
  assign _T_1057 = reset | io_reset;
  assign _T_1064 = ~ SRFF_io_output_data;
  assign _T_1065 = ~ denseLoadBuffers_0_io_deqVld;
  assign _T_1074 = denseLoadBuffers_0_io_deqVld & _T_1068;
  assign _T_1075 = _T_1064 & _T_1074;
  assign _T_1079 = ~ SRFF_1_io_output_data;
  assign _T_1080 = ~ denseLoadBuffers_0_io_enqVld;
  assign _T_1089 = denseLoadBuffers_0_io_enqVld & _T_1083;
  assign _T_1090 = _T_1079 & _T_1089;
  assign _T_1091 = {denseLoadBuffers_0_io_enq_15,denseLoadBuffers_0_io_enq_14};
  assign _T_1092 = {_T_1091,denseLoadBuffers_0_io_enq_13};
  assign _T_1093 = {_T_1092,denseLoadBuffers_0_io_enq_12};
  assign _T_1094 = {_T_1093,denseLoadBuffers_0_io_enq_11};
  assign _T_1095 = {_T_1094,denseLoadBuffers_0_io_enq_10};
  assign _T_1096 = {_T_1095,denseLoadBuffers_0_io_enq_9};
  assign _T_1097 = {_T_1096,denseLoadBuffers_0_io_enq_8};
  assign _T_1098 = {_T_1097,denseLoadBuffers_0_io_enq_7};
  assign _T_1099 = {_T_1098,denseLoadBuffers_0_io_enq_6};
  assign _T_1100 = {_T_1099,denseLoadBuffers_0_io_enq_5};
  assign _T_1101 = {_T_1100,denseLoadBuffers_0_io_enq_4};
  assign _T_1102 = {_T_1101,denseLoadBuffers_0_io_enq_3};
  assign _T_1103 = {_T_1102,denseLoadBuffers_0_io_enq_2};
  assign _T_1104 = {_T_1103,denseLoadBuffers_0_io_enq_1};
  assign _T_1105 = {_T_1104,denseLoadBuffers_0_io_enq_0};
  assign _T_1109 = burstCounterDoneLatch_io_out & sizeCounterDoneLatch_io_out;
  assign _T_1110 = cmdWrite & wdataMux_io_out_valid;
  assign _T_1111 = ~ dramReadySeen;
  assign _T_1112 = _T_1110 & _T_1111;
  assign _T_1114 = ~ denseStoreBuffers_0_io_empty;
  assign _T_1115 = cmdWrite & _T_1114;
  assign _T_1116 = _T_1115 & io_dram_wdata_ready;
  assign _T_1118 = cmdArbiter_io_tag;
  assign _T_1119 = _T_1116 & _T_1118;
  assign _T_1120 = ~ cmdCooldown_io_out;
  assign _T_1121 = _T_1119 & _T_1120;
  assign _T_1122 = ~ burstCounterDoneLatch_io_out;
  assign _T_1123 = _T_1121 & _T_1122;
  assign _T_1127 = _T_1115 & _T_1120;
  assign _T_1129 = _T_1127 & _T_1122;
  assign _T_1130 = denseStoreBuffers_0_io_deqStrb[0];
  assign _T_1131 = denseStoreBuffers_0_io_deqStrb[1];
  assign _T_1132 = denseStoreBuffers_0_io_deqStrb[2];
  assign _T_1133 = denseStoreBuffers_0_io_deqStrb[3];
  assign _T_1134 = denseStoreBuffers_0_io_deqStrb[4];
  assign _T_1135 = denseStoreBuffers_0_io_deqStrb[5];
  assign _T_1136 = denseStoreBuffers_0_io_deqStrb[6];
  assign _T_1137 = denseStoreBuffers_0_io_deqStrb[7];
  assign _T_1138 = denseStoreBuffers_0_io_deqStrb[8];
  assign _T_1139 = denseStoreBuffers_0_io_deqStrb[9];
  assign _T_1140 = denseStoreBuffers_0_io_deqStrb[10];
  assign _T_1141 = denseStoreBuffers_0_io_deqStrb[11];
  assign _T_1142 = denseStoreBuffers_0_io_deqStrb[12];
  assign _T_1143 = denseStoreBuffers_0_io_deqStrb[13];
  assign _T_1144 = denseStoreBuffers_0_io_deqStrb[14];
  assign _T_1145 = denseStoreBuffers_0_io_deqStrb[15];
  assign _T_1146 = denseStoreBuffers_0_io_deqStrb[16];
  assign _T_1147 = denseStoreBuffers_0_io_deqStrb[17];
  assign _T_1148 = denseStoreBuffers_0_io_deqStrb[18];
  assign _T_1149 = denseStoreBuffers_0_io_deqStrb[19];
  assign _T_1150 = denseStoreBuffers_0_io_deqStrb[20];
  assign _T_1151 = denseStoreBuffers_0_io_deqStrb[21];
  assign _T_1152 = denseStoreBuffers_0_io_deqStrb[22];
  assign _T_1153 = denseStoreBuffers_0_io_deqStrb[23];
  assign _T_1154 = denseStoreBuffers_0_io_deqStrb[24];
  assign _T_1155 = denseStoreBuffers_0_io_deqStrb[25];
  assign _T_1156 = denseStoreBuffers_0_io_deqStrb[26];
  assign _T_1157 = denseStoreBuffers_0_io_deqStrb[27];
  assign _T_1158 = denseStoreBuffers_0_io_deqStrb[28];
  assign _T_1159 = denseStoreBuffers_0_io_deqStrb[29];
  assign _T_1160 = denseStoreBuffers_0_io_deqStrb[30];
  assign _T_1161 = denseStoreBuffers_0_io_deqStrb[31];
  assign _T_1162 = denseStoreBuffers_0_io_deqStrb[32];
  assign _T_1163 = denseStoreBuffers_0_io_deqStrb[33];
  assign _T_1164 = denseStoreBuffers_0_io_deqStrb[34];
  assign _T_1165 = denseStoreBuffers_0_io_deqStrb[35];
  assign _T_1166 = denseStoreBuffers_0_io_deqStrb[36];
  assign _T_1167 = denseStoreBuffers_0_io_deqStrb[37];
  assign _T_1168 = denseStoreBuffers_0_io_deqStrb[38];
  assign _T_1169 = denseStoreBuffers_0_io_deqStrb[39];
  assign _T_1170 = denseStoreBuffers_0_io_deqStrb[40];
  assign _T_1171 = denseStoreBuffers_0_io_deqStrb[41];
  assign _T_1172 = denseStoreBuffers_0_io_deqStrb[42];
  assign _T_1173 = denseStoreBuffers_0_io_deqStrb[43];
  assign _T_1174 = denseStoreBuffers_0_io_deqStrb[44];
  assign _T_1175 = denseStoreBuffers_0_io_deqStrb[45];
  assign _T_1176 = denseStoreBuffers_0_io_deqStrb[46];
  assign _T_1177 = denseStoreBuffers_0_io_deqStrb[47];
  assign _T_1178 = denseStoreBuffers_0_io_deqStrb[48];
  assign _T_1179 = denseStoreBuffers_0_io_deqStrb[49];
  assign _T_1180 = denseStoreBuffers_0_io_deqStrb[50];
  assign _T_1181 = denseStoreBuffers_0_io_deqStrb[51];
  assign _T_1182 = denseStoreBuffers_0_io_deqStrb[52];
  assign _T_1183 = denseStoreBuffers_0_io_deqStrb[53];
  assign _T_1184 = denseStoreBuffers_0_io_deqStrb[54];
  assign _T_1185 = denseStoreBuffers_0_io_deqStrb[55];
  assign _T_1186 = denseStoreBuffers_0_io_deqStrb[56];
  assign _T_1187 = denseStoreBuffers_0_io_deqStrb[57];
  assign _T_1188 = denseStoreBuffers_0_io_deqStrb[58];
  assign _T_1189 = denseStoreBuffers_0_io_deqStrb[59];
  assign _T_1190 = denseStoreBuffers_0_io_deqStrb[60];
  assign _T_1191 = denseStoreBuffers_0_io_deqStrb[61];
  assign _T_1192 = denseStoreBuffers_0_io_deqStrb[62];
  assign _T_1193 = denseStoreBuffers_0_io_deqStrb[63];
  assign _T_1194 = ~ denseStoreBuffers_0_io_full;
  assign _T_1197 = io_dram_cmd_valid & io_dram_cmd_ready;
  assign _T_1202 = io_dram_wresp_bits_tag_streamId == 6'h1;
  assign _T_1203 = io_dram_wresp_valid & _T_1202;
  assign _T_1204 = ~ FIFOCounter_io_full;
  assign _T_1205 = ~ FIFOCounter_io_empty;
  assign burstCounterMax = _T_1197 ? io_dram_cmd_bits_size : burstCounterMaxLatch_io_out;
  assign _T_1227 = isSparseMux_io_out ? 1'h0 : burstCounter_io_done;
  assign _T_1229 = burstCounter_io_last ? _T_1109 : burstCounterDoneLatch_io_out;
  assign _T_1231 = io_dram_cmd_bits_isWr ? burstCounterMax : 32'h1;
  assign _T_1233 = wdataMux_io_out_valid & io_dram_wdata_ready;
  assign _T_1235 = io_dram_cmd_bits_isWr ? _T_1233 : _T_1197;
  assign dramReadyFFEnabler = isSparseMux_io_out ? burstCounter_io_done : burstCounterDoneLatch_io_out;
  assign _T_1243 = io_dram_cmd_valid & io_dram_cmd_bits_isWr;
  assign _T_1244 = dramReadyFFEnabler | _T_1243;
  assign _T_1246 = io_dram_cmd_ready | dramReadySeen;
  assign _T_1247 = dramReadyFFEnabler ? 1'h0 : _T_1246;
  assign _T_1249 = ~ _T_1197;
  assign _T_1255 = isSparseMux_io_out ? 1'h1 : _T_1120;
  assign _T_1256 = dramCmdMux_io_out_valid & _T_1255;
  assign _T_1261 = io_dram_rresp_valid & io_dram_rresp_ready;
  assign _T_1266 = io_dram_wdata_valid & io_dram_wdata_ready;
  assign _T_1267 = _T_1266 & io_enable;
  assign _T_1272 = io_enable & io_dram_cmd_ready;
  assign _T_1273 = _T_1272 & io_dram_cmd_valid;
  assign _T_1278 = ~ cmdArbiter_io_empty;
  assign _T_1279 = io_enable & _T_1278;
  assign _T_1280 = io_dram_cmd_ready & io_dram_cmd_valid;
  assign _T_1281 = ~ _T_1280;
  assign _T_1282 = _T_1279 & _T_1281;
  assign _T_1290 = _T_1273 & _T_897;
  assign _T_1295 = io_enable & io_app_loads_0_cmd_valid;
  assign _T_1301 = _T_1295 & io_app_loads_0_cmd_ready;
  assign _T_1308 = cmdArbiter_io_tag == 1'h0;
  assign _T_1309 = _T_1197 & _T_1308;
  assign _T_1316 = _T_1273 & cmdArbiter_io_deq_0_isWr;
  assign _T_1335 = _T_1197 & _T_1118;
  assign _T_1345 = io_enable & io_dram_rresp_valid;
  assign _T_1346 = ~ io_dram_rresp_ready;
  assign _T_1347 = _T_1345 & _T_1346;
  assign _T_1352 = ~ io_dram_rresp_valid;
  assign _T_1353 = io_enable & _T_1352;
  assign _T_1354 = _T_1353 & io_dram_rresp_ready;
  assign _T_1362 = _T_1261 & _T_1027;
  assign _T_1367 = io_dram_wresp_valid & io_dram_wresp_ready;
  assign _T_1372 = io_enable & io_dram_wresp_valid;
  assign _T_1373 = ~ io_dram_wresp_ready;
  assign _T_1374 = _T_1372 & _T_1373;
  assign _T_1379 = ~ io_dram_wresp_valid;
  assign _T_1380 = io_enable & _T_1379;
  assign _T_1381 = _T_1380 & io_dram_wresp_ready;
  assign _T_1389 = _T_1367 & _T_1202;
  assign _T_1425 = io_dram_rresp_bits_tag_streamId >= 6'h1;
  assign _T_1443 = _T_1194 & denseStoreBuffers_0_io_enqVld;
  assign _T_1448 = denseStoreBuffers_0_io_full & denseStoreBuffers_0_io_enqVld;
  assign _T_1469 = io_dram_rresp_valid & denseLoadBuffers_0_io_enqVld;
  assign _T_1480 = _T_1261 & denseLoadBuffers_0_io_enqVld;
  assign _T_1486 = io_dram_rresp_valid & _T_1346;
  assign io_app_loads_0_cmd_ready = _T_891;
  assign io_app_loads_0_rdata_valid = _T_1031;
  assign io_app_loads_0_rdata_bits_0 = denseLoadBuffers_0_io_deq_0;
  assign io_dram_cmd_valid = _T_1256;
  assign io_dram_cmd_bits_addr = dramCmdMux_io_out_bits_addr;
  assign io_dram_cmd_bits_size = dramCmdMux_io_out_bits_size;
  assign io_dram_cmd_bits_isWr = dramCmdMux_io_out_bits_isWr;
  assign io_dram_cmd_bits_tag_uid = dramCmdMux_io_out_bits_tag_uid;
  assign io_dram_cmd_bits_tag_streamId = dramCmdMux_io_out_bits_tag_streamId;
  assign io_dram_wdata_valid = wdataMux_io_out_valid;
  assign io_dram_wdata_bits_wdata_0 = wdataMux_io_out_bits_wdata_0;
  assign io_dram_wdata_bits_wdata_1 = wdataMux_io_out_bits_wdata_1;
  assign io_dram_wdata_bits_wdata_2 = wdataMux_io_out_bits_wdata_2;
  assign io_dram_wdata_bits_wdata_3 = wdataMux_io_out_bits_wdata_3;
  assign io_dram_wdata_bits_wdata_4 = wdataMux_io_out_bits_wdata_4;
  assign io_dram_wdata_bits_wdata_5 = wdataMux_io_out_bits_wdata_5;
  assign io_dram_wdata_bits_wdata_6 = wdataMux_io_out_bits_wdata_6;
  assign io_dram_wdata_bits_wdata_7 = wdataMux_io_out_bits_wdata_7;
  assign io_dram_wdata_bits_wdata_8 = wdataMux_io_out_bits_wdata_8;
  assign io_dram_wdata_bits_wdata_9 = wdataMux_io_out_bits_wdata_9;
  assign io_dram_wdata_bits_wdata_10 = wdataMux_io_out_bits_wdata_10;
  assign io_dram_wdata_bits_wdata_11 = wdataMux_io_out_bits_wdata_11;
  assign io_dram_wdata_bits_wdata_12 = wdataMux_io_out_bits_wdata_12;
  assign io_dram_wdata_bits_wdata_13 = wdataMux_io_out_bits_wdata_13;
  assign io_dram_wdata_bits_wdata_14 = wdataMux_io_out_bits_wdata_14;
  assign io_dram_wdata_bits_wdata_15 = wdataMux_io_out_bits_wdata_15;
  assign io_dram_wdata_bits_wstrb_0 = wdataMux_io_out_bits_wstrb_63;
  assign io_dram_wdata_bits_wstrb_1 = wdataMux_io_out_bits_wstrb_62;
  assign io_dram_wdata_bits_wstrb_2 = wdataMux_io_out_bits_wstrb_61;
  assign io_dram_wdata_bits_wstrb_3 = wdataMux_io_out_bits_wstrb_60;
  assign io_dram_wdata_bits_wstrb_4 = wdataMux_io_out_bits_wstrb_59;
  assign io_dram_wdata_bits_wstrb_5 = wdataMux_io_out_bits_wstrb_58;
  assign io_dram_wdata_bits_wstrb_6 = wdataMux_io_out_bits_wstrb_57;
  assign io_dram_wdata_bits_wstrb_7 = wdataMux_io_out_bits_wstrb_56;
  assign io_dram_wdata_bits_wstrb_8 = wdataMux_io_out_bits_wstrb_55;
  assign io_dram_wdata_bits_wstrb_9 = wdataMux_io_out_bits_wstrb_54;
  assign io_dram_wdata_bits_wstrb_10 = wdataMux_io_out_bits_wstrb_53;
  assign io_dram_wdata_bits_wstrb_11 = wdataMux_io_out_bits_wstrb_52;
  assign io_dram_wdata_bits_wstrb_12 = wdataMux_io_out_bits_wstrb_51;
  assign io_dram_wdata_bits_wstrb_13 = wdataMux_io_out_bits_wstrb_50;
  assign io_dram_wdata_bits_wstrb_14 = wdataMux_io_out_bits_wstrb_49;
  assign io_dram_wdata_bits_wstrb_15 = wdataMux_io_out_bits_wstrb_48;
  assign io_dram_wdata_bits_wstrb_16 = wdataMux_io_out_bits_wstrb_47;
  assign io_dram_wdata_bits_wstrb_17 = wdataMux_io_out_bits_wstrb_46;
  assign io_dram_wdata_bits_wstrb_18 = wdataMux_io_out_bits_wstrb_45;
  assign io_dram_wdata_bits_wstrb_19 = wdataMux_io_out_bits_wstrb_44;
  assign io_dram_wdata_bits_wstrb_20 = wdataMux_io_out_bits_wstrb_43;
  assign io_dram_wdata_bits_wstrb_21 = wdataMux_io_out_bits_wstrb_42;
  assign io_dram_wdata_bits_wstrb_22 = wdataMux_io_out_bits_wstrb_41;
  assign io_dram_wdata_bits_wstrb_23 = wdataMux_io_out_bits_wstrb_40;
  assign io_dram_wdata_bits_wstrb_24 = wdataMux_io_out_bits_wstrb_39;
  assign io_dram_wdata_bits_wstrb_25 = wdataMux_io_out_bits_wstrb_38;
  assign io_dram_wdata_bits_wstrb_26 = wdataMux_io_out_bits_wstrb_37;
  assign io_dram_wdata_bits_wstrb_27 = wdataMux_io_out_bits_wstrb_36;
  assign io_dram_wdata_bits_wstrb_28 = wdataMux_io_out_bits_wstrb_35;
  assign io_dram_wdata_bits_wstrb_29 = wdataMux_io_out_bits_wstrb_34;
  assign io_dram_wdata_bits_wstrb_30 = wdataMux_io_out_bits_wstrb_33;
  assign io_dram_wdata_bits_wstrb_31 = wdataMux_io_out_bits_wstrb_32;
  assign io_dram_wdata_bits_wstrb_32 = wdataMux_io_out_bits_wstrb_31;
  assign io_dram_wdata_bits_wstrb_33 = wdataMux_io_out_bits_wstrb_30;
  assign io_dram_wdata_bits_wstrb_34 = wdataMux_io_out_bits_wstrb_29;
  assign io_dram_wdata_bits_wstrb_35 = wdataMux_io_out_bits_wstrb_28;
  assign io_dram_wdata_bits_wstrb_36 = wdataMux_io_out_bits_wstrb_27;
  assign io_dram_wdata_bits_wstrb_37 = wdataMux_io_out_bits_wstrb_26;
  assign io_dram_wdata_bits_wstrb_38 = wdataMux_io_out_bits_wstrb_25;
  assign io_dram_wdata_bits_wstrb_39 = wdataMux_io_out_bits_wstrb_24;
  assign io_dram_wdata_bits_wstrb_40 = wdataMux_io_out_bits_wstrb_23;
  assign io_dram_wdata_bits_wstrb_41 = wdataMux_io_out_bits_wstrb_22;
  assign io_dram_wdata_bits_wstrb_42 = wdataMux_io_out_bits_wstrb_21;
  assign io_dram_wdata_bits_wstrb_43 = wdataMux_io_out_bits_wstrb_20;
  assign io_dram_wdata_bits_wstrb_44 = wdataMux_io_out_bits_wstrb_19;
  assign io_dram_wdata_bits_wstrb_45 = wdataMux_io_out_bits_wstrb_18;
  assign io_dram_wdata_bits_wstrb_46 = wdataMux_io_out_bits_wstrb_17;
  assign io_dram_wdata_bits_wstrb_47 = wdataMux_io_out_bits_wstrb_16;
  assign io_dram_wdata_bits_wstrb_48 = wdataMux_io_out_bits_wstrb_15;
  assign io_dram_wdata_bits_wstrb_49 = wdataMux_io_out_bits_wstrb_14;
  assign io_dram_wdata_bits_wstrb_50 = wdataMux_io_out_bits_wstrb_13;
  assign io_dram_wdata_bits_wstrb_51 = wdataMux_io_out_bits_wstrb_12;
  assign io_dram_wdata_bits_wstrb_52 = wdataMux_io_out_bits_wstrb_11;
  assign io_dram_wdata_bits_wstrb_53 = wdataMux_io_out_bits_wstrb_10;
  assign io_dram_wdata_bits_wstrb_54 = wdataMux_io_out_bits_wstrb_9;
  assign io_dram_wdata_bits_wstrb_55 = wdataMux_io_out_bits_wstrb_8;
  assign io_dram_wdata_bits_wstrb_56 = wdataMux_io_out_bits_wstrb_7;
  assign io_dram_wdata_bits_wstrb_57 = wdataMux_io_out_bits_wstrb_6;
  assign io_dram_wdata_bits_wstrb_58 = wdataMux_io_out_bits_wstrb_5;
  assign io_dram_wdata_bits_wstrb_59 = wdataMux_io_out_bits_wstrb_4;
  assign io_dram_wdata_bits_wstrb_60 = wdataMux_io_out_bits_wstrb_3;
  assign io_dram_wdata_bits_wstrb_61 = wdataMux_io_out_bits_wstrb_2;
  assign io_dram_wdata_bits_wstrb_62 = wdataMux_io_out_bits_wstrb_1;
  assign io_dram_wdata_bits_wstrb_63 = wdataMux_io_out_bits_wstrb_0;
  assign io_dram_rresp_ready = rrespReadyMux_io_out;
  assign io_dram_wresp_ready = wrespReadyMux_io_out;
  assign cmdArbiter_io_fifo_0_deq_0_addr = cmdFifos_0_io_deq_0_addr;
  assign cmdArbiter_io_fifo_0_deq_0_isWr = cmdFifos_0_io_deq_0_isWr;
  assign cmdArbiter_io_fifo_0_deq_0_size = cmdFifos_0_io_deq_0_size;
  assign cmdArbiter_io_fifo_0_full = cmdFifos_0_io_full;
  assign cmdArbiter_io_fifo_0_empty = cmdFifos_0_io_empty;
  assign cmdArbiter_io_fifo_0_almostEmpty = cmdFifos_0_io_almostEmpty;
  assign cmdArbiter_io_fifo_1_deq_0_addr = cmdFifos_1_io_deq_0_addr;
  assign cmdArbiter_io_fifo_1_deq_0_isWr = cmdFifos_1_io_deq_0_isWr;
  assign cmdArbiter_io_fifo_1_deq_0_size = cmdFifos_1_io_deq_0_size;
  assign cmdArbiter_io_fifo_1_empty = cmdFifos_1_io_empty;
  assign cmdArbiter_io_enq_0_0_addr = io_app_loads_0_cmd_bits_addr;
  assign cmdArbiter_io_enq_0_0_isWr = io_app_loads_0_cmd_bits_isWr;
  assign cmdArbiter_io_enq_0_0_size = io_app_loads_0_cmd_bits_size;
  assign cmdArbiter_io_enqVld_0 = io_app_loads_0_cmd_valid;
  assign cmdArbiter_io_deqVld = cmdDeqValidMux_io_out;
  assign cmdArbiter_clock = clock;
  assign cmdArbiter_reset = reset;
  assign cmdFifos_0_io_enq_0_addr = cmdArbiter_io_fifo_0_enq_0_addr;
  assign cmdFifos_0_io_enq_0_isWr = cmdArbiter_io_fifo_0_enq_0_isWr;
  assign cmdFifos_0_io_enq_0_size = cmdArbiter_io_fifo_0_enq_0_size;
  assign cmdFifos_0_io_enqVld = cmdArbiter_io_fifo_0_enqVld;
  assign cmdFifos_0_io_deqVld = cmdArbiter_io_fifo_0_deqVld;
  assign cmdFifos_0_clock = clock;
  assign cmdFifos_0_reset = reset;
  assign cmdFifos_1_io_enq_0_addr = 64'h0;
  assign cmdFifos_1_io_enq_0_isWr = 1'h0;
  assign cmdFifos_1_io_enq_0_size = 16'h0;
  assign cmdFifos_1_io_enqVld = 1'h0;
  assign cmdFifos_1_io_deqVld = cmdArbiter_io_fifo_1_deqVld;
  assign cmdFifos_1_clock = clock;
  assign cmdFifos_1_reset = reset;
  assign FF_io_in = _T_887;
  assign FF_io_init = 64'h175be;
  assign FF_io_reset = 1'h0;
  assign FF_io_enable = io_app_loads_0_cmd_valid;
  assign FF_clock = clock;
  assign FF_reset = reset;
  assign sizeCounter_io_max = _T_903;
  assign sizeCounter_io_stride = 16'h4000;
  assign sizeCounter_io_reset = 1'h0;
  assign sizeCounter_io_enable = _T_1197;
  assign sizeCounter_clock = clock;
  assign sizeCounter_reset = reset;
  assign cmdAddr_bits = _T_895;
  assign isSparseMux_io_ins_0 = 1'h0;
  assign isSparseMux_io_ins_1 = 1'h0;
  assign isSparseMux_io_sel = cmdArbiter_io_tag;
  assign burstCounter_io_max = _T_1231[15:0];
  assign burstCounter_io_stride = 16'h1;
  assign burstCounter_io_reset = io_reset;
  assign burstCounter_io_enable = _T_1235;
  assign burstCounter_clock = clock;
  assign burstCounter_reset = reset;
  assign burstTagCounter_io_reset = io_reset;
  assign burstTagCounter_io_enable = _T_1197;
  assign burstTagCounter_clock = clock;
  assign burstTagCounter_reset = reset;
  assign dramReadySeen = dramReadyFF_io_out;
  assign cmdCooldown_io_in = 1'h1;
  assign cmdCooldown_io_init = 1'h0;
  assign cmdCooldown_io_reset = _T_1249;
  assign cmdCooldown_io_enable = _T_1197;
  assign cmdCooldown_clock = clock;
  assign cmdCooldown_reset = reset;
  assign burstCounterDoneLatch_io_in = 1'h1;
  assign burstCounterDoneLatch_io_init = 1'h0;
  assign burstCounterDoneLatch_io_reset = _T_1229;
  assign burstCounterDoneLatch_io_enable = _T_1227;
  assign burstCounterDoneLatch_clock = clock;
  assign burstCounterDoneLatch_reset = reset;
  assign sizeCounterDoneLatch_io_in = 1'h1;
  assign sizeCounterDoneLatch_io_init = 1'h0;
  assign sizeCounterDoneLatch_io_reset = burstCounterDoneLatch_io_out;
  assign sizeCounterDoneLatch_io_enable = _T_908;
  assign sizeCounterDoneLatch_clock = clock;
  assign sizeCounterDoneLatch_reset = reset;
  assign rrespReadyMux_io_ins_0 = _T_1029;
  assign wdataMux_io_ins_0_valid = _T_1129;
  assign wdataMux_io_ins_0_bits_wdata_0 = denseStoreBuffers_0_io_deq_0;
  assign wdataMux_io_ins_0_bits_wdata_1 = denseStoreBuffers_0_io_deq_1;
  assign wdataMux_io_ins_0_bits_wdata_2 = denseStoreBuffers_0_io_deq_2;
  assign wdataMux_io_ins_0_bits_wdata_3 = denseStoreBuffers_0_io_deq_3;
  assign wdataMux_io_ins_0_bits_wdata_4 = denseStoreBuffers_0_io_deq_4;
  assign wdataMux_io_ins_0_bits_wdata_5 = denseStoreBuffers_0_io_deq_5;
  assign wdataMux_io_ins_0_bits_wdata_6 = denseStoreBuffers_0_io_deq_6;
  assign wdataMux_io_ins_0_bits_wdata_7 = denseStoreBuffers_0_io_deq_7;
  assign wdataMux_io_ins_0_bits_wdata_8 = denseStoreBuffers_0_io_deq_8;
  assign wdataMux_io_ins_0_bits_wdata_9 = denseStoreBuffers_0_io_deq_9;
  assign wdataMux_io_ins_0_bits_wdata_10 = denseStoreBuffers_0_io_deq_10;
  assign wdataMux_io_ins_0_bits_wdata_11 = denseStoreBuffers_0_io_deq_11;
  assign wdataMux_io_ins_0_bits_wdata_12 = denseStoreBuffers_0_io_deq_12;
  assign wdataMux_io_ins_0_bits_wdata_13 = denseStoreBuffers_0_io_deq_13;
  assign wdataMux_io_ins_0_bits_wdata_14 = denseStoreBuffers_0_io_deq_14;
  assign wdataMux_io_ins_0_bits_wdata_15 = denseStoreBuffers_0_io_deq_15;
  assign wdataMux_io_ins_0_bits_wstrb_0 = _T_1130;
  assign wdataMux_io_ins_0_bits_wstrb_1 = _T_1131;
  assign wdataMux_io_ins_0_bits_wstrb_2 = _T_1132;
  assign wdataMux_io_ins_0_bits_wstrb_3 = _T_1133;
  assign wdataMux_io_ins_0_bits_wstrb_4 = _T_1134;
  assign wdataMux_io_ins_0_bits_wstrb_5 = _T_1135;
  assign wdataMux_io_ins_0_bits_wstrb_6 = _T_1136;
  assign wdataMux_io_ins_0_bits_wstrb_7 = _T_1137;
  assign wdataMux_io_ins_0_bits_wstrb_8 = _T_1138;
  assign wdataMux_io_ins_0_bits_wstrb_9 = _T_1139;
  assign wdataMux_io_ins_0_bits_wstrb_10 = _T_1140;
  assign wdataMux_io_ins_0_bits_wstrb_11 = _T_1141;
  assign wdataMux_io_ins_0_bits_wstrb_12 = _T_1142;
  assign wdataMux_io_ins_0_bits_wstrb_13 = _T_1143;
  assign wdataMux_io_ins_0_bits_wstrb_14 = _T_1144;
  assign wdataMux_io_ins_0_bits_wstrb_15 = _T_1145;
  assign wdataMux_io_ins_0_bits_wstrb_16 = _T_1146;
  assign wdataMux_io_ins_0_bits_wstrb_17 = _T_1147;
  assign wdataMux_io_ins_0_bits_wstrb_18 = _T_1148;
  assign wdataMux_io_ins_0_bits_wstrb_19 = _T_1149;
  assign wdataMux_io_ins_0_bits_wstrb_20 = _T_1150;
  assign wdataMux_io_ins_0_bits_wstrb_21 = _T_1151;
  assign wdataMux_io_ins_0_bits_wstrb_22 = _T_1152;
  assign wdataMux_io_ins_0_bits_wstrb_23 = _T_1153;
  assign wdataMux_io_ins_0_bits_wstrb_24 = _T_1154;
  assign wdataMux_io_ins_0_bits_wstrb_25 = _T_1155;
  assign wdataMux_io_ins_0_bits_wstrb_26 = _T_1156;
  assign wdataMux_io_ins_0_bits_wstrb_27 = _T_1157;
  assign wdataMux_io_ins_0_bits_wstrb_28 = _T_1158;
  assign wdataMux_io_ins_0_bits_wstrb_29 = _T_1159;
  assign wdataMux_io_ins_0_bits_wstrb_30 = _T_1160;
  assign wdataMux_io_ins_0_bits_wstrb_31 = _T_1161;
  assign wdataMux_io_ins_0_bits_wstrb_32 = _T_1162;
  assign wdataMux_io_ins_0_bits_wstrb_33 = _T_1163;
  assign wdataMux_io_ins_0_bits_wstrb_34 = _T_1164;
  assign wdataMux_io_ins_0_bits_wstrb_35 = _T_1165;
  assign wdataMux_io_ins_0_bits_wstrb_36 = _T_1166;
  assign wdataMux_io_ins_0_bits_wstrb_37 = _T_1167;
  assign wdataMux_io_ins_0_bits_wstrb_38 = _T_1168;
  assign wdataMux_io_ins_0_bits_wstrb_39 = _T_1169;
  assign wdataMux_io_ins_0_bits_wstrb_40 = _T_1170;
  assign wdataMux_io_ins_0_bits_wstrb_41 = _T_1171;
  assign wdataMux_io_ins_0_bits_wstrb_42 = _T_1172;
  assign wdataMux_io_ins_0_bits_wstrb_43 = _T_1173;
  assign wdataMux_io_ins_0_bits_wstrb_44 = _T_1174;
  assign wdataMux_io_ins_0_bits_wstrb_45 = _T_1175;
  assign wdataMux_io_ins_0_bits_wstrb_46 = _T_1176;
  assign wdataMux_io_ins_0_bits_wstrb_47 = _T_1177;
  assign wdataMux_io_ins_0_bits_wstrb_48 = _T_1178;
  assign wdataMux_io_ins_0_bits_wstrb_49 = _T_1179;
  assign wdataMux_io_ins_0_bits_wstrb_50 = _T_1180;
  assign wdataMux_io_ins_0_bits_wstrb_51 = _T_1181;
  assign wdataMux_io_ins_0_bits_wstrb_52 = _T_1182;
  assign wdataMux_io_ins_0_bits_wstrb_53 = _T_1183;
  assign wdataMux_io_ins_0_bits_wstrb_54 = _T_1184;
  assign wdataMux_io_ins_0_bits_wstrb_55 = _T_1185;
  assign wdataMux_io_ins_0_bits_wstrb_56 = _T_1186;
  assign wdataMux_io_ins_0_bits_wstrb_57 = _T_1187;
  assign wdataMux_io_ins_0_bits_wstrb_58 = _T_1188;
  assign wdataMux_io_ins_0_bits_wstrb_59 = _T_1189;
  assign wdataMux_io_ins_0_bits_wstrb_60 = _T_1190;
  assign wdataMux_io_ins_0_bits_wstrb_61 = _T_1191;
  assign wdataMux_io_ins_0_bits_wstrb_62 = _T_1192;
  assign wdataMux_io_ins_0_bits_wstrb_63 = _T_1193;
  assign cmdDeqValidMux_io_ins_0 = sizeCounterDoneLatch_io_out;
  assign cmdDeqValidMux_io_ins_1 = _T_1109;
  assign cmdDeqValidMux_io_sel = cmdArbiter_io_tag;
  assign dramCmdMux_io_ins_0_valid = cmdRead;
  assign dramCmdMux_io_ins_0_bits_addr = _T_933;
  assign dramCmdMux_io_ins_0_bits_size = {{22'd0}, _T_949};
  assign dramCmdMux_io_ins_0_bits_isWr = cmdArbiter_io_deq_0_isWr;
  assign dramCmdMux_io_ins_0_bits_tag_uid = {{16'd0}, burstTagCounter_io_out};
  assign dramCmdMux_io_ins_0_bits_tag_streamId = _T_935_streamId;
  assign dramCmdMux_io_ins_1_valid = _T_1112;
  assign dramCmdMux_io_ins_1_bits_addr = _T_933;
  assign dramCmdMux_io_ins_1_bits_size = {{22'd0}, _T_983};
  assign dramCmdMux_io_ins_1_bits_isWr = cmdArbiter_io_deq_0_isWr;
  assign dramCmdMux_io_ins_1_bits_tag_uid = {{16'd0}, burstTagCounter_io_out};
  assign dramCmdMux_io_ins_1_bits_tag_streamId = _T_969_streamId;
  assign dramCmdMux_io_sel = cmdArbiter_io_tag;
  assign _T_935_streamId = {{5'd0}, cmdArbiter_io_tag};
  assign _T_937_bits = _T_943;
  assign FF_1_io_in = dramCmdMux_io_out_bits_tag_streamId;
  assign FF_1_io_enable = _T_951;
  assign FF_1_clock = clock;
  assign FF_1_reset = reset;
  assign FF_2_io_in = dramCmdMux_io_out_bits_addr;
  assign FF_2_io_init = 64'h175be;
  assign FF_2_io_reset = 1'h0;
  assign FF_2_io_enable = _T_951;
  assign FF_2_clock = clock;
  assign FF_2_reset = reset;
  assign FF_3_io_in = dramCmdMux_io_out_bits_size;
  assign FF_3_io_enable = _T_951;
  assign FF_3_clock = clock;
  assign FF_3_reset = reset;
  assign _T_969_streamId = {{5'd0}, cmdArbiter_io_tag};
  assign _T_971_bits = _T_943;
  assign FF_4_io_in = cmdArbiter_io_tag;
  assign FF_4_io_init = 1'h0;
  assign FF_4_io_reset = 1'h0;
  assign FF_4_io_enable = cmdWrite;
  assign FF_4_clock = clock;
  assign FF_4_reset = reset;
  assign FF_5_io_in = cmdArbiter_io_deq_0_size;
  assign FF_5_io_enable = cmdWrite;
  assign FF_5_clock = clock;
  assign FF_5_reset = reset;
  assign wrespReadyMux_io_ins_0 = _T_1204;
  assign gatherLoadIssueMux_io_ins_0 = 1'h0;
  assign gatherLoadIssueMux_io_ins_1 = 1'h0;
  assign gatherLoadIssueMux_io_sel = cmdArbiter_io_tag;
  assign gatherLoadIssue_io_reset = io_reset;
  assign gatherLoadIssue_io_enable = gatherLoadIssueMux_io_out;
  assign gatherLoadIssue_clock = clock;
  assign gatherLoadIssue_reset = reset;
  assign gatherLoadSkipMux_io_ins_0 = 1'h0;
  assign gatherLoadSkipMux_io_ins_1 = 1'h0;
  assign gatherLoadSkipMux_io_sel = cmdArbiter_io_tag;
  assign gatherLoadSkip_io_reset = io_reset;
  assign gatherLoadSkip_io_enable = gatherLoadSkipMux_io_out;
  assign gatherLoadSkip_clock = clock;
  assign gatherLoadSkip_reset = reset;
  assign scatterLoadIssueMux_io_ins_0 = 1'h0;
  assign scatterLoadIssueMux_io_ins_1 = 1'h0;
  assign scatterLoadIssueMux_io_sel = cmdArbiter_io_tag;
  assign scatterLoadIssue_io_reset = io_reset;
  assign scatterLoadIssue_io_enable = scatterLoadIssueMux_io_out;
  assign scatterLoadIssue_clock = clock;
  assign scatterLoadIssue_reset = reset;
  assign scatterLoadSkipMux_io_ins_0 = 1'h0;
  assign scatterLoadSkipMux_io_ins_1 = 1'h0;
  assign scatterLoadSkipMux_io_sel = cmdArbiter_io_tag;
  assign scatterLoadSkip_io_reset = io_reset;
  assign scatterLoadSkip_io_enable = scatterLoadSkipMux_io_out;
  assign scatterLoadSkip_clock = clock;
  assign scatterLoadSkip_reset = reset;
  assign scatterStoreIssueMux_io_ins_0 = 1'h0;
  assign scatterStoreIssueMux_io_ins_1 = 1'h0;
  assign scatterStoreIssueMux_io_sel = cmdArbiter_io_tag;
  assign scatterStoreIssue_io_reset = io_reset;
  assign scatterStoreIssue_io_enable = scatterStoreIssueMux_io_out;
  assign scatterStoreIssue_clock = clock;
  assign scatterStoreIssue_reset = reset;
  assign scatterStoreSkipMux_io_ins_0 = 1'h0;
  assign scatterStoreSkipMux_io_ins_1 = 1'h0;
  assign scatterStoreSkipMux_io_sel = cmdArbiter_io_tag;
  assign scatterStoreSkip_io_reset = io_reset;
  assign scatterStoreSkip_io_enable = scatterStoreSkipMux_io_out;
  assign scatterStoreSkip_clock = clock;
  assign scatterStoreSkip_reset = reset;
  assign denseLoadBuffers_0_io_enq_0 = io_dram_rresp_bits_rdata_0;
  assign denseLoadBuffers_0_io_enq_1 = io_dram_rresp_bits_rdata_1;
  assign denseLoadBuffers_0_io_enq_2 = io_dram_rresp_bits_rdata_2;
  assign denseLoadBuffers_0_io_enq_3 = io_dram_rresp_bits_rdata_3;
  assign denseLoadBuffers_0_io_enq_4 = io_dram_rresp_bits_rdata_4;
  assign denseLoadBuffers_0_io_enq_5 = io_dram_rresp_bits_rdata_5;
  assign denseLoadBuffers_0_io_enq_6 = io_dram_rresp_bits_rdata_6;
  assign denseLoadBuffers_0_io_enq_7 = io_dram_rresp_bits_rdata_7;
  assign denseLoadBuffers_0_io_enq_8 = io_dram_rresp_bits_rdata_8;
  assign denseLoadBuffers_0_io_enq_9 = io_dram_rresp_bits_rdata_9;
  assign denseLoadBuffers_0_io_enq_10 = io_dram_rresp_bits_rdata_10;
  assign denseLoadBuffers_0_io_enq_11 = io_dram_rresp_bits_rdata_11;
  assign denseLoadBuffers_0_io_enq_12 = io_dram_rresp_bits_rdata_12;
  assign denseLoadBuffers_0_io_enq_13 = io_dram_rresp_bits_rdata_13;
  assign denseLoadBuffers_0_io_enq_14 = io_dram_rresp_bits_rdata_14;
  assign denseLoadBuffers_0_io_enq_15 = io_dram_rresp_bits_rdata_15;
  assign denseLoadBuffers_0_io_enqVld = _T_1028;
  assign denseLoadBuffers_0_io_deqVld = io_app_loads_0_rdata_ready;
  assign denseLoadBuffers_0_clock = clock;
  assign denseLoadBuffers_0_reset = reset;
  assign Counter_io_reset = io_reset;
  assign Counter_io_enable = denseLoadBuffers_0_io_enqVld;
  assign Counter_clock = clock;
  assign Counter_reset = reset;
  assign Counter_1_io_reset = io_reset;
  assign Counter_1_io_enable = _T_1031;
  assign Counter_1_clock = clock;
  assign Counter_1_reset = reset;
  assign Counter_2_io_reset = io_reset;
  assign Counter_2_io_enable = io_app_loads_0_rdata_ready;
  assign Counter_2_clock = clock;
  assign Counter_2_reset = reset;
  assign Counter_3_io_reset = io_reset;
  assign Counter_3_io_enable = _T_1046;
  assign Counter_3_clock = clock;
  assign Counter_3_reset = reset;
  assign Counter_4_io_reset = io_reset;
  assign Counter_4_io_enable = _T_1051;
  assign Counter_4_clock = clock;
  assign Counter_4_reset = reset;
  assign SRFF_io_input_set = denseLoadBuffers_0_io_deqVld;
  assign SRFF_io_input_reset = _T_1057;
  assign SRFF_io_input_asyn_reset = _T_1057;
  assign SRFF_clock = clock;
  assign SRFF_reset = reset;
  assign SRFF_1_io_input_set = denseLoadBuffers_0_io_enqVld;
  assign SRFF_1_io_input_reset = _T_1057;
  assign SRFF_1_io_input_asyn_reset = _T_1057;
  assign SRFF_1_clock = clock;
  assign SRFF_1_reset = reset;
  assign FF_6_io_in = denseLoadBuffers_0_io_deq_0;
  assign FF_6_io_enable = _T_1075;
  assign FF_6_clock = clock;
  assign FF_6_reset = reset;
  assign FF_7_io_in = _T_1105;
  assign FF_7_io_enable = _T_1090;
  assign FF_7_clock = clock;
  assign FF_7_reset = reset;
  assign denseStoreBuffers_0_io_enqVld = 1'h0;
  assign denseStoreBuffers_0_io_deqVld = _T_1123;
  assign denseStoreBuffers_0_clock = clock;
  assign denseStoreBuffers_0_reset = reset;
  assign Counter_5_io_max = FF_8_io_out;
  assign Counter_5_io_stride = 16'h4000;
  assign Counter_5_io_reset = 1'h0;
  assign Counter_5_io_enable = _T_1203;
  assign Counter_5_clock = clock;
  assign Counter_5_reset = reset;
  assign FF_8_io_in = cmdArbiter_io_deq_0_size;
  assign FF_8_io_enable = _T_1197;
  assign FF_8_clock = clock;
  assign FF_8_reset = reset;
  assign FIFOCounter_io_enqVld = Counter_5_io_done;
  assign FIFOCounter_clock = clock;
  assign FIFOCounter_reset = reset;
  assign Counter_6_io_reset = io_reset;
  assign Counter_6_io_enable = FIFOCounter_io_enqVld;
  assign Counter_6_clock = clock;
  assign Counter_6_reset = reset;
  assign Counter_7_io_reset = io_reset;
  assign Counter_7_io_enable = _T_1205;
  assign Counter_7_clock = clock;
  assign Counter_7_reset = reset;
  assign Counter_8_io_reset = io_reset;
  assign Counter_8_io_enable = 1'h0;
  assign Counter_8_clock = clock;
  assign Counter_8_reset = reset;
  assign burstCounterMaxLatch_io_in = io_dram_cmd_bits_size;
  assign burstCounterMaxLatch_io_enable = _T_1197;
  assign burstCounterMaxLatch_clock = clock;
  assign burstCounterMaxLatch_reset = reset;
  assign dramReadyFF_io_in = _T_1247;
  assign dramReadyFF_io_init = 1'h0;
  assign dramReadyFF_io_reset = 1'h0;
  assign dramReadyFF_io_enable = _T_1244;
  assign dramReadyFF_clock = clock;
  assign dramReadyFF_reset = reset;
  assign cycleCount_io_reset = io_reset;
  assign cycleCount_io_enable = io_enable;
  assign cycleCount_clock = clock;
  assign cycleCount_reset = reset;
  assign rdataEnqCount_io_reset = io_reset;
  assign rdataEnqCount_io_enable = _T_1261;
  assign rdataEnqCount_clock = clock;
  assign rdataEnqCount_reset = reset;
  assign wdataCount_io_reset = io_reset;
  assign wdataCount_io_enable = _T_1267;
  assign wdataCount_clock = clock;
  assign wdataCount_reset = reset;
  assign Counter_9_io_reset = io_reset;
  assign Counter_9_io_enable = _T_1273;
  assign Counter_9_clock = clock;
  assign Counter_9_reset = reset;
  assign Counter_10_io_reset = io_reset;
  assign Counter_10_io_enable = _T_1282;
  assign Counter_10_clock = clock;
  assign Counter_10_reset = reset;
  assign Counter_11_io_reset = io_reset;
  assign Counter_11_io_enable = _T_1290;
  assign Counter_11_clock = clock;
  assign Counter_11_reset = reset;
  assign Counter_12_io_reset = io_reset;
  assign Counter_12_io_enable = _T_1295;
  assign Counter_12_clock = clock;
  assign Counter_12_reset = reset;
  assign Counter_13_io_reset = io_reset;
  assign Counter_13_io_enable = _T_1301;
  assign Counter_13_clock = clock;
  assign Counter_13_reset = reset;
  assign Counter_14_io_reset = io_reset;
  assign Counter_14_io_enable = _T_1309;
  assign Counter_14_clock = clock;
  assign Counter_14_reset = reset;
  assign Counter_15_io_reset = io_reset;
  assign Counter_15_io_enable = _T_1316;
  assign Counter_15_clock = clock;
  assign Counter_15_reset = reset;
  assign Counter_16_io_reset = io_reset;
  assign Counter_16_io_enable = 1'h0;
  assign Counter_16_clock = clock;
  assign Counter_16_reset = reset;
  assign Counter_17_io_reset = io_reset;
  assign Counter_17_io_enable = 1'h0;
  assign Counter_17_clock = clock;
  assign Counter_17_reset = reset;
  assign Counter_18_io_reset = io_reset;
  assign Counter_18_io_enable = _T_1335;
  assign Counter_18_clock = clock;
  assign Counter_18_reset = reset;
  assign Counter_19_io_reset = io_reset;
  assign Counter_19_io_enable = _T_1261;
  assign Counter_19_clock = clock;
  assign Counter_19_reset = reset;
  assign Counter_20_io_reset = io_reset;
  assign Counter_20_io_enable = _T_1347;
  assign Counter_20_clock = clock;
  assign Counter_20_reset = reset;
  assign Counter_21_io_reset = io_reset;
  assign Counter_21_io_enable = _T_1354;
  assign Counter_21_clock = clock;
  assign Counter_21_reset = reset;
  assign Counter_22_io_reset = io_reset;
  assign Counter_22_io_enable = _T_1362;
  assign Counter_22_clock = clock;
  assign Counter_22_reset = reset;
  assign Counter_23_io_reset = io_reset;
  assign Counter_23_io_enable = _T_1367;
  assign Counter_23_clock = clock;
  assign Counter_23_reset = reset;
  assign Counter_24_io_reset = io_reset;
  assign Counter_24_io_enable = _T_1374;
  assign Counter_24_clock = clock;
  assign Counter_24_reset = reset;
  assign Counter_25_io_reset = io_reset;
  assign Counter_25_io_enable = _T_1381;
  assign Counter_25_clock = clock;
  assign Counter_25_reset = reset;
  assign Counter_26_io_reset = io_reset;
  assign Counter_26_io_enable = _T_1389;
  assign Counter_26_clock = clock;
  assign Counter_26_reset = reset;
  assign Counter_27_io_reset = io_reset;
  assign Counter_27_io_enable = denseLoadBuffers_0_io_full;
  assign Counter_27_clock = clock;
  assign Counter_27_reset = reset;
  assign Counter_28_io_reset = io_reset;
  assign Counter_28_io_enable = denseLoadBuffers_0_io_almostFull;
  assign Counter_28_clock = clock;
  assign Counter_28_reset = reset;
  assign Counter_29_io_reset = io_reset;
  assign Counter_29_io_enable = denseLoadBuffers_0_io_empty;
  assign Counter_29_clock = clock;
  assign Counter_29_reset = reset;
  assign Counter_30_io_reset = io_reset;
  assign Counter_30_io_enable = denseLoadBuffers_0_io_almostEmpty;
  assign Counter_30_clock = clock;
  assign Counter_30_reset = reset;
  assign Counter_31_io_reset = io_reset;
  assign Counter_31_io_enable = denseLoadBuffers_0_io_enqVld;
  assign Counter_31_clock = clock;
  assign Counter_31_reset = reset;
  assign Counter_32_io_reset = io_reset;
  assign Counter_32_io_enable = _T_1027;
  assign Counter_32_clock = clock;
  assign Counter_32_reset = reset;
  assign Counter_33_io_reset = io_reset;
  assign Counter_33_io_enable = io_dram_rresp_valid;
  assign Counter_33_clock = clock;
  assign Counter_33_reset = reset;
  assign Counter_34_io_reset = io_reset;
  assign Counter_34_io_enable = _T_1425;
  assign Counter_34_clock = clock;
  assign Counter_34_reset = reset;
  assign FF_9_io_in = io_dram_rresp_bits_tag_streamId;
  assign FF_9_io_enable = io_dram_rresp_valid;
  assign FF_9_clock = clock;
  assign FF_9_reset = reset;
  assign Counter_35_io_reset = io_reset;
  assign Counter_35_io_enable = denseStoreBuffers_0_io_enqVld;
  assign Counter_35_clock = clock;
  assign Counter_35_reset = reset;
  assign Counter_36_io_reset = io_reset;
  assign Counter_36_io_enable = _T_1194;
  assign Counter_36_clock = clock;
  assign Counter_36_reset = reset;
  assign Counter_37_io_reset = io_reset;
  assign Counter_37_io_enable = _T_1443;
  assign Counter_37_clock = clock;
  assign Counter_37_reset = reset;
  assign Counter_38_io_reset = io_reset;
  assign Counter_38_io_enable = _T_1448;
  assign Counter_38_clock = clock;
  assign Counter_38_reset = reset;
  assign Counter_39_io_reset = io_reset;
  assign Counter_39_io_enable = denseStoreBuffers_0_io_full;
  assign Counter_39_clock = clock;
  assign Counter_39_reset = reset;
  assign Counter_40_io_reset = io_reset;
  assign Counter_40_io_enable = denseStoreBuffers_0_io_almostFull;
  assign Counter_40_clock = clock;
  assign Counter_40_reset = reset;
  assign Counter_41_io_reset = io_reset;
  assign Counter_41_io_enable = denseStoreBuffers_0_io_empty;
  assign Counter_41_clock = clock;
  assign Counter_41_reset = reset;
  assign Counter_42_io_reset = io_reset;
  assign Counter_42_io_enable = denseStoreBuffers_0_io_almostEmpty;
  assign Counter_42_clock = clock;
  assign Counter_42_reset = reset;
  assign Counter_43_io_reset = io_reset;
  assign Counter_43_io_enable = _T_1469;
  assign Counter_43_clock = clock;
  assign Counter_43_reset = reset;
  assign Counter_44_io_reset = io_reset;
  assign Counter_44_io_enable = _T_1261;
  assign Counter_44_clock = clock;
  assign Counter_44_reset = reset;
  assign Counter_45_io_reset = io_reset;
  assign Counter_45_io_enable = _T_1480;
  assign Counter_45_clock = clock;
  assign Counter_45_reset = reset;
  assign Counter_46_io_reset = io_reset;
  assign Counter_46_io_enable = _T_1486;
  assign Counter_46_clock = clock;
  assign Counter_46_reset = reset;
  assign Counter_47_io_reset = io_reset;
  assign Counter_47_io_enable = 1'h0;
  assign Counter_47_clock = clock;
  assign Counter_47_reset = reset;
  assign Counter_48_io_reset = io_reset;
  assign Counter_48_io_enable = 1'h0;
  assign Counter_48_clock = clock;
  assign Counter_48_reset = reset;
  assign Counter_49_io_reset = io_reset;
  assign Counter_49_io_enable = 1'h0;
  assign Counter_49_clock = clock;
  assign Counter_49_reset = reset;
  assign Counter_50_io_reset = io_reset;
  assign Counter_50_io_enable = 1'h0;
  assign Counter_50_clock = clock;
  assign Counter_50_reset = reset;
  assign Counter_51_io_reset = io_reset;
  assign Counter_51_io_enable = 1'h0;
  assign Counter_51_clock = clock;
  assign Counter_51_reset = reset;
  assign Counter_52_io_reset = io_reset;
  assign Counter_52_io_enable = 1'h0;
  assign Counter_52_clock = clock;
  assign Counter_52_reset = reset;
  assign Counter_53_io_reset = io_reset;
  assign Counter_53_io_enable = 1'h0;
  assign Counter_53_clock = clock;
  assign Counter_53_reset = reset;
  assign Counter_54_io_reset = io_reset;
  assign Counter_54_io_enable = 1'h0;
  assign Counter_54_clock = clock;
  assign Counter_54_reset = reset;
  assign Counter_55_io_reset = io_reset;
  assign Counter_55_io_enable = 1'h0;
  assign Counter_55_clock = clock;
  assign Counter_55_reset = reset;
  assign Counter_56_io_reset = io_reset;
  assign Counter_56_io_enable = 1'h0;
  assign Counter_56_clock = clock;
  assign Counter_56_reset = reset;
  assign Counter_57_io_reset = io_reset;
  assign Counter_57_io_enable = 1'h1;
  assign Counter_57_clock = clock;
  assign Counter_57_reset = reset;
  assign Counter_58_io_reset = io_reset;
  assign Counter_58_io_enable = 1'h0;
  assign Counter_58_clock = clock;
  assign Counter_58_reset = reset;
  assign Counter_59_io_reset = io_reset;
  assign Counter_59_io_enable = 1'h0;
  assign Counter_59_clock = clock;
  assign Counter_59_reset = reset;
  assign FF_10_io_in = 64'h0;
  assign FF_10_io_init = 64'h175be;
  assign FF_10_io_reset = 1'h0;
  assign FF_10_io_enable = 1'h0;
  assign FF_10_clock = clock;
  assign FF_10_reset = reset;
  assign FF_11_io_in = 8'h0;
  assign FF_11_io_enable = 1'h0;
  assign FF_11_clock = clock;
  assign FF_11_reset = reset;
  assign FF_12_io_in = 3'h0;
  assign FF_12_io_enable = 1'h0;
  assign FF_12_clock = clock;
  assign FF_12_reset = reset;
  assign FF_13_io_in = 1'h0;
  assign FF_13_io_init = 1'h0;
  assign FF_13_io_reset = 1'h0;
  assign FF_13_io_enable = 1'h0;
  assign FF_13_clock = clock;
  assign FF_13_reset = reset;
  assign FF_14_io_in = 2'h0;
  assign FF_14_io_enable = 1'h0;
  assign FF_14_clock = clock;
  assign FF_14_reset = reset;
  assign FF_15_io_in = 64'h0;
  assign FF_15_io_init = 64'h175be;
  assign FF_15_io_reset = 1'h0;
  assign FF_15_io_enable = 1'h0;
  assign FF_15_clock = clock;
  assign FF_15_reset = reset;
  assign FF_16_io_in = 8'h0;
  assign FF_16_io_enable = 1'h0;
  assign FF_16_clock = clock;
  assign FF_16_reset = reset;
  assign FF_17_io_in = 512'h0;
  assign FF_17_io_enable = 1'h0;
  assign FF_17_clock = clock;
  assign FF_17_reset = reset;
  assign FF_18_io_in = 64'h0;
  assign FF_18_io_init = 64'h175be;
  assign FF_18_io_reset = 1'h0;
  assign FF_18_io_enable = 1'h0;
  assign FF_18_clock = clock;
  assign FF_18_reset = reset;
  assign FF_19_io_in = 512'h0;
  assign FF_19_io_enable = 1'h0;
  assign FF_19_clock = clock;
  assign FF_19_reset = reset;
  assign FF_20_io_in = 64'h0;
  assign FF_20_io_init = 64'h175be;
  assign FF_20_io_reset = 1'h0;
  assign FF_20_io_enable = 1'h0;
  assign FF_20_clock = clock;
  assign FF_20_reset = reset;
  assign FF_21_io_in = 512'h0;
  assign FF_21_io_enable = 1'h0;
  assign FF_21_clock = clock;
  assign FF_21_reset = reset;
  assign FF_22_io_in = 64'h0;
  assign FF_22_io_init = 64'h175be;
  assign FF_22_io_reset = 1'h0;
  assign FF_22_io_enable = 1'h0;
  assign FF_22_clock = clock;
  assign FF_22_reset = reset;
  assign Counter_60_io_reset = io_reset;
  assign Counter_60_io_enable = 1'h0;
  assign Counter_60_clock = clock;
  assign Counter_60_reset = reset;
  assign Counter_61_io_reset = io_reset;
  assign Counter_61_io_enable = 1'h0;
  assign Counter_61_clock = clock;
  assign Counter_61_reset = reset;
  assign Counter_62_io_reset = io_reset;
  assign Counter_62_io_enable = 1'h0;
  assign Counter_62_clock = clock;
  assign Counter_62_reset = reset;
  assign Counter_63_io_reset = io_reset;
  assign Counter_63_io_enable = 1'h0;
  assign Counter_63_clock = clock;
  assign Counter_63_reset = reset;
  assign Counter_64_io_reset = io_reset;
  assign Counter_64_io_enable = 1'h0;
  assign Counter_64_clock = clock;
  assign Counter_64_reset = reset;
  assign Counter_65_io_reset = io_reset;
  assign Counter_65_io_enable = 1'h0;
  assign Counter_65_clock = clock;
  assign Counter_65_reset = reset;
  assign Counter_66_io_reset = io_reset;
  assign Counter_66_io_enable = 1'h0;
  assign Counter_66_clock = clock;
  assign Counter_66_reset = reset;
  assign Counter_67_io_reset = io_reset;
  assign Counter_67_io_enable = 1'h0;
  assign Counter_67_clock = clock;
  assign Counter_67_reset = reset;
  assign Counter_68_io_reset = io_reset;
  assign Counter_68_io_enable = 1'h0;
  assign Counter_68_clock = clock;
  assign Counter_68_reset = reset;
  assign Counter_69_io_reset = io_reset;
  assign Counter_69_io_enable = 1'h0;
  assign Counter_69_clock = clock;
  assign Counter_69_reset = reset;
  assign Counter_70_io_reset = io_reset;
  assign Counter_70_io_enable = 1'h1;
  assign Counter_70_clock = clock;
  assign Counter_70_reset = reset;
  assign Counter_71_io_reset = io_reset;
  assign Counter_71_io_enable = 1'h0;
  assign Counter_71_clock = clock;
  assign Counter_71_reset = reset;
  assign Counter_72_io_reset = io_reset;
  assign Counter_72_io_enable = 1'h0;
  assign Counter_72_clock = clock;
  assign Counter_72_reset = reset;
  assign FF_23_io_in = 64'h0;
  assign FF_23_io_init = 64'h175be;
  assign FF_23_io_reset = 1'h0;
  assign FF_23_io_enable = 1'h0;
  assign FF_23_clock = clock;
  assign FF_23_reset = reset;
  assign FF_24_io_in = 8'h0;
  assign FF_24_io_enable = 1'h0;
  assign FF_24_clock = clock;
  assign FF_24_reset = reset;
  assign FF_25_io_in = 3'h0;
  assign FF_25_io_enable = 1'h0;
  assign FF_25_clock = clock;
  assign FF_25_reset = reset;
  assign FF_26_io_in = 2'h0;
  assign FF_26_io_enable = 1'h0;
  assign FF_26_clock = clock;
  assign FF_26_reset = reset;
  assign FF_27_io_in = 64'h0;
  assign FF_27_io_init = 64'h175be;
  assign FF_27_io_reset = 1'h0;
  assign FF_27_io_enable = 1'h0;
  assign FF_27_clock = clock;
  assign FF_27_reset = reset;
  assign FF_28_io_in = 8'h0;
  assign FF_28_io_enable = 1'h0;
  assign FF_28_clock = clock;
  assign FF_28_reset = reset;
  assign FF_29_io_in = 512'h0;
  assign FF_29_io_enable = 1'h0;
  assign FF_29_clock = clock;
  assign FF_29_reset = reset;
  assign FF_30_io_in = 64'h0;
  assign FF_30_io_init = 64'h175be;
  assign FF_30_io_reset = 1'h0;
  assign FF_30_io_enable = 1'h0;
  assign FF_30_clock = clock;
  assign FF_30_reset = reset;
  assign FF_31_io_in = 512'h0;
  assign FF_31_io_enable = 1'h0;
  assign FF_31_clock = clock;
  assign FF_31_reset = reset;
  assign FF_32_io_in = 64'h0;
  assign FF_32_io_init = 64'h175be;
  assign FF_32_io_reset = 1'h0;
  assign FF_32_io_enable = 1'h0;
  assign FF_32_clock = clock;
  assign FF_32_reset = reset;
  assign FF_33_io_in = 512'h0;
  assign FF_33_io_enable = 1'h0;
  assign FF_33_clock = clock;
  assign FF_33_reset = reset;
  assign FF_34_io_in = 64'h0;
  assign FF_34_io_init = 64'h175be;
  assign FF_34_io_reset = 1'h0;
  assign FF_34_io_enable = 1'h0;
  assign FF_34_clock = clock;
  assign FF_34_reset = reset;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_1068 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_1083 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_1068 <= 1'h0;
    end else begin
      _T_1068 <= _T_1065;
    end
    if (reset) begin
      _T_1083 <= 1'h0;
    end else begin
      _T_1083 <= _T_1080;
    end
  end
endmodule
module MuxN_80(
  input  [63:0] io_ins_0,
  input  [63:0] io_ins_1,
  input  [63:0] io_ins_2,
  input  [63:0] io_ins_3,
  input  [63:0] io_ins_4,
  input  [63:0] io_ins_5,
  input  [63:0] io_ins_6,
  input  [63:0] io_ins_7,
  input  [63:0] io_ins_8,
  input  [63:0] io_ins_9,
  input  [63:0] io_ins_10,
  input  [63:0] io_ins_11,
  input  [63:0] io_ins_12,
  input  [63:0] io_ins_13,
  input  [63:0] io_ins_14,
  input  [63:0] io_ins_15,
  input  [63:0] io_ins_16,
  input  [63:0] io_ins_17,
  input  [63:0] io_ins_18,
  input  [63:0] io_ins_19,
  input  [63:0] io_ins_20,
  input  [63:0] io_ins_21,
  input  [63:0] io_ins_22,
  input  [63:0] io_ins_23,
  input  [63:0] io_ins_24,
  input  [63:0] io_ins_25,
  input  [63:0] io_ins_26,
  input  [63:0] io_ins_27,
  input  [63:0] io_ins_28,
  input  [63:0] io_ins_29,
  input  [63:0] io_ins_30,
  input  [63:0] io_ins_31,
  input  [63:0] io_ins_32,
  input  [63:0] io_ins_33,
  input  [63:0] io_ins_34,
  input  [63:0] io_ins_35,
  input  [63:0] io_ins_36,
  input  [63:0] io_ins_37,
  input  [63:0] io_ins_38,
  input  [63:0] io_ins_39,
  input  [63:0] io_ins_40,
  input  [63:0] io_ins_41,
  input  [63:0] io_ins_42,
  input  [63:0] io_ins_43,
  input  [63:0] io_ins_44,
  input  [63:0] io_ins_45,
  input  [63:0] io_ins_46,
  input  [63:0] io_ins_47,
  input  [63:0] io_ins_48,
  input  [63:0] io_ins_49,
  input  [63:0] io_ins_50,
  input  [63:0] io_ins_51,
  input  [63:0] io_ins_52,
  input  [63:0] io_ins_53,
  input  [63:0] io_ins_54,
  input  [63:0] io_ins_55,
  input  [63:0] io_ins_56,
  input  [63:0] io_ins_57,
  input  [63:0] io_ins_58,
  input  [63:0] io_ins_59,
  input  [63:0] io_ins_60,
  input  [63:0] io_ins_61,
  input  [63:0] io_ins_62,
  input  [63:0] io_ins_63,
  input  [63:0] io_ins_64,
  input  [63:0] io_ins_65,
  input  [63:0] io_ins_66,
  input  [63:0] io_ins_67,
  input  [63:0] io_ins_68,
  input  [63:0] io_ins_69,
  input  [63:0] io_ins_70,
  input  [63:0] io_ins_71,
  input  [63:0] io_ins_72,
  input  [63:0] io_ins_73,
  input  [63:0] io_ins_74,
  input  [63:0] io_ins_75,
  input  [63:0] io_ins_76,
  input  [63:0] io_ins_77,
  input  [63:0] io_ins_78,
  input  [63:0] io_ins_79,
  input  [63:0] io_ins_80,
  input  [63:0] io_ins_81,
  input  [63:0] io_ins_82,
  input  [63:0] io_ins_83,
  input  [63:0] io_ins_84,
  input  [63:0] io_ins_85,
  input  [63:0] io_ins_86,
  input  [63:0] io_ins_87,
  input  [63:0] io_ins_88,
  input  [63:0] io_ins_89,
  input  [63:0] io_ins_90,
  input  [63:0] io_ins_91,
  input  [63:0] io_ins_92,
  input  [63:0] io_ins_93,
  input  [63:0] io_ins_94,
  input  [63:0] io_ins_95,
  input  [63:0] io_ins_96,
  input  [63:0] io_ins_97,
  input  [63:0] io_ins_98,
  input  [63:0] io_ins_99,
  input  [63:0] io_ins_100,
  input  [63:0] io_ins_101,
  input  [63:0] io_ins_102,
  input  [63:0] io_ins_103,
  input  [63:0] io_ins_104,
  input  [63:0] io_ins_105,
  input  [63:0] io_ins_106,
  input  [63:0] io_ins_107,
  input  [63:0] io_ins_108,
  input  [63:0] io_ins_109,
  input  [63:0] io_ins_110,
  input  [63:0] io_ins_111,
  input  [63:0] io_ins_112,
  input  [63:0] io_ins_113,
  input  [63:0] io_ins_114,
  input  [63:0] io_ins_115,
  input  [63:0] io_ins_116,
  input  [63:0] io_ins_117,
  input  [63:0] io_ins_118,
  input  [63:0] io_ins_119,
  input  [63:0] io_ins_120,
  input  [63:0] io_ins_121,
  input  [63:0] io_ins_122,
  input  [63:0] io_ins_123,
  input  [63:0] io_ins_124,
  input  [63:0] io_ins_125,
  input  [63:0] io_ins_126,
  input  [63:0] io_ins_127,
  input  [63:0] io_ins_128,
  input  [63:0] io_ins_129,
  input  [63:0] io_ins_130,
  input  [63:0] io_ins_131,
  input  [63:0] io_ins_132,
  input  [63:0] io_ins_133,
  input  [63:0] io_ins_134,
  input  [63:0] io_ins_135,
  input  [63:0] io_ins_136,
  input  [63:0] io_ins_137,
  input  [63:0] io_ins_138,
  input  [63:0] io_ins_139,
  input  [63:0] io_ins_140,
  input  [63:0] io_ins_141,
  input  [63:0] io_ins_142,
  input  [63:0] io_ins_143,
  input  [63:0] io_ins_144,
  input  [63:0] io_ins_145,
  input  [63:0] io_ins_146,
  input  [63:0] io_ins_147,
  input  [63:0] io_ins_148,
  input  [63:0] io_ins_149,
  input  [63:0] io_ins_150,
  input  [63:0] io_ins_151,
  input  [63:0] io_ins_152,
  input  [63:0] io_ins_153,
  input  [63:0] io_ins_154,
  input  [63:0] io_ins_155,
  input  [63:0] io_ins_156,
  input  [63:0] io_ins_157,
  input  [63:0] io_ins_158,
  input  [63:0] io_ins_159,
  input  [63:0] io_ins_160,
  input  [63:0] io_ins_161,
  input  [63:0] io_ins_162,
  input  [63:0] io_ins_163,
  input  [63:0] io_ins_164,
  input  [63:0] io_ins_165,
  input  [63:0] io_ins_166,
  input  [63:0] io_ins_167,
  input  [63:0] io_ins_168,
  input  [63:0] io_ins_169,
  input  [63:0] io_ins_170,
  input  [63:0] io_ins_171,
  input  [63:0] io_ins_172,
  input  [63:0] io_ins_173,
  input  [63:0] io_ins_174,
  input  [63:0] io_ins_175,
  input  [63:0] io_ins_176,
  input  [63:0] io_ins_177,
  input  [63:0] io_ins_178,
  input  [63:0] io_ins_179,
  input  [63:0] io_ins_180,
  input  [63:0] io_ins_181,
  input  [63:0] io_ins_182,
  input  [63:0] io_ins_183,
  input  [63:0] io_ins_184,
  input  [63:0] io_ins_185,
  input  [63:0] io_ins_186,
  input  [63:0] io_ins_187,
  input  [63:0] io_ins_188,
  input  [63:0] io_ins_189,
  input  [63:0] io_ins_190,
  input  [63:0] io_ins_191,
  input  [63:0] io_ins_192,
  input  [63:0] io_ins_193,
  input  [63:0] io_ins_194,
  input  [63:0] io_ins_195,
  input  [63:0] io_ins_196,
  input  [63:0] io_ins_197,
  input  [63:0] io_ins_198,
  input  [63:0] io_ins_199,
  input  [63:0] io_ins_200,
  input  [63:0] io_ins_201,
  input  [63:0] io_ins_202,
  input  [63:0] io_ins_203,
  input  [63:0] io_ins_204,
  input  [63:0] io_ins_205,
  input  [63:0] io_ins_206,
  input  [63:0] io_ins_207,
  input  [63:0] io_ins_208,
  input  [63:0] io_ins_209,
  input  [63:0] io_ins_210,
  input  [63:0] io_ins_211,
  input  [63:0] io_ins_212,
  input  [63:0] io_ins_213,
  input  [63:0] io_ins_214,
  input  [63:0] io_ins_215,
  input  [63:0] io_ins_216,
  input  [63:0] io_ins_217,
  input  [63:0] io_ins_218,
  input  [63:0] io_ins_219,
  input  [63:0] io_ins_220,
  input  [63:0] io_ins_221,
  input  [63:0] io_ins_222,
  input  [63:0] io_ins_223,
  input  [63:0] io_ins_224,
  input  [63:0] io_ins_225,
  input  [63:0] io_ins_226,
  input  [63:0] io_ins_227,
  input  [63:0] io_ins_228,
  input  [63:0] io_ins_229,
  input  [63:0] io_ins_230,
  input  [63:0] io_ins_231,
  input  [63:0] io_ins_232,
  input  [63:0] io_ins_233,
  input  [63:0] io_ins_234,
  input  [63:0] io_ins_235,
  input  [63:0] io_ins_236,
  input  [63:0] io_ins_237,
  input  [63:0] io_ins_238,
  input  [63:0] io_ins_239,
  input  [63:0] io_ins_240,
  input  [63:0] io_ins_241,
  input  [63:0] io_ins_242,
  input  [63:0] io_ins_243,
  input  [63:0] io_ins_244,
  input  [63:0] io_ins_245,
  input  [63:0] io_ins_246,
  input  [63:0] io_ins_247,
  input  [63:0] io_ins_248,
  input  [63:0] io_ins_249,
  input  [63:0] io_ins_250,
  input  [63:0] io_ins_251,
  input  [63:0] io_ins_252,
  input  [63:0] io_ins_253,
  input  [63:0] io_ins_254,
  input  [63:0] io_ins_255,
  input  [63:0] io_ins_256,
  input  [63:0] io_ins_257,
  input  [63:0] io_ins_258,
  input  [63:0] io_ins_259,
  input  [63:0] io_ins_260,
  input  [63:0] io_ins_261,
  input  [63:0] io_ins_262,
  input  [63:0] io_ins_263,
  input  [63:0] io_ins_264,
  input  [63:0] io_ins_265,
  input  [63:0] io_ins_266,
  input  [63:0] io_ins_267,
  input  [63:0] io_ins_268,
  input  [63:0] io_ins_269,
  input  [63:0] io_ins_270,
  input  [63:0] io_ins_271,
  input  [63:0] io_ins_272,
  input  [63:0] io_ins_273,
  input  [63:0] io_ins_274,
  input  [63:0] io_ins_275,
  input  [63:0] io_ins_276,
  input  [63:0] io_ins_277,
  input  [63:0] io_ins_278,
  input  [63:0] io_ins_279,
  input  [63:0] io_ins_280,
  input  [63:0] io_ins_281,
  input  [63:0] io_ins_282,
  input  [63:0] io_ins_283,
  input  [63:0] io_ins_284,
  input  [63:0] io_ins_285,
  input  [63:0] io_ins_286,
  input  [63:0] io_ins_287,
  input  [63:0] io_ins_288,
  input  [63:0] io_ins_289,
  input  [63:0] io_ins_290,
  input  [63:0] io_ins_291,
  input  [63:0] io_ins_292,
  input  [63:0] io_ins_293,
  input  [63:0] io_ins_294,
  input  [63:0] io_ins_295,
  input  [63:0] io_ins_296,
  input  [63:0] io_ins_297,
  input  [63:0] io_ins_298,
  input  [63:0] io_ins_299,
  input  [63:0] io_ins_300,
  input  [63:0] io_ins_301,
  input  [63:0] io_ins_302,
  input  [63:0] io_ins_303,
  input  [63:0] io_ins_304,
  input  [63:0] io_ins_305,
  input  [63:0] io_ins_306,
  input  [63:0] io_ins_307,
  input  [63:0] io_ins_308,
  input  [63:0] io_ins_309,
  input  [63:0] io_ins_310,
  input  [63:0] io_ins_311,
  input  [63:0] io_ins_312,
  input  [63:0] io_ins_313,
  input  [63:0] io_ins_314,
  input  [63:0] io_ins_315,
  input  [63:0] io_ins_316,
  input  [63:0] io_ins_317,
  input  [63:0] io_ins_318,
  input  [63:0] io_ins_319,
  input  [63:0] io_ins_320,
  input  [63:0] io_ins_321,
  input  [63:0] io_ins_322,
  input  [63:0] io_ins_323,
  input  [63:0] io_ins_324,
  input  [63:0] io_ins_325,
  input  [63:0] io_ins_326,
  input  [63:0] io_ins_327,
  input  [63:0] io_ins_328,
  input  [63:0] io_ins_329,
  input  [63:0] io_ins_330,
  input  [63:0] io_ins_331,
  input  [63:0] io_ins_332,
  input  [63:0] io_ins_333,
  input  [63:0] io_ins_334,
  input  [63:0] io_ins_335,
  input  [63:0] io_ins_336,
  input  [63:0] io_ins_337,
  input  [63:0] io_ins_338,
  input  [63:0] io_ins_339,
  input  [63:0] io_ins_340,
  input  [63:0] io_ins_341,
  input  [63:0] io_ins_342,
  input  [63:0] io_ins_343,
  input  [63:0] io_ins_344,
  input  [63:0] io_ins_345,
  input  [63:0] io_ins_346,
  input  [63:0] io_ins_347,
  input  [63:0] io_ins_348,
  input  [63:0] io_ins_349,
  input  [63:0] io_ins_350,
  input  [63:0] io_ins_351,
  input  [63:0] io_ins_352,
  input  [63:0] io_ins_353,
  input  [63:0] io_ins_354,
  input  [63:0] io_ins_355,
  input  [63:0] io_ins_356,
  input  [63:0] io_ins_357,
  input  [63:0] io_ins_358,
  input  [63:0] io_ins_359,
  input  [63:0] io_ins_360,
  input  [63:0] io_ins_361,
  input  [63:0] io_ins_362,
  input  [63:0] io_ins_363,
  input  [63:0] io_ins_364,
  input  [63:0] io_ins_365,
  input  [63:0] io_ins_366,
  input  [63:0] io_ins_367,
  input  [63:0] io_ins_368,
  input  [63:0] io_ins_369,
  input  [63:0] io_ins_370,
  input  [63:0] io_ins_371,
  input  [63:0] io_ins_372,
  input  [63:0] io_ins_373,
  input  [63:0] io_ins_374,
  input  [63:0] io_ins_375,
  input  [63:0] io_ins_376,
  input  [63:0] io_ins_377,
  input  [63:0] io_ins_378,
  input  [63:0] io_ins_379,
  input  [63:0] io_ins_380,
  input  [63:0] io_ins_381,
  input  [63:0] io_ins_382,
  input  [63:0] io_ins_383,
  input  [63:0] io_ins_384,
  input  [63:0] io_ins_385,
  input  [63:0] io_ins_386,
  input  [63:0] io_ins_387,
  input  [63:0] io_ins_388,
  input  [63:0] io_ins_389,
  input  [63:0] io_ins_390,
  input  [63:0] io_ins_391,
  input  [63:0] io_ins_392,
  input  [63:0] io_ins_393,
  input  [63:0] io_ins_394,
  input  [63:0] io_ins_395,
  input  [63:0] io_ins_396,
  input  [63:0] io_ins_397,
  input  [63:0] io_ins_398,
  input  [63:0] io_ins_399,
  input  [63:0] io_ins_400,
  input  [63:0] io_ins_401,
  input  [63:0] io_ins_402,
  input  [63:0] io_ins_403,
  input  [63:0] io_ins_404,
  input  [63:0] io_ins_405,
  input  [63:0] io_ins_406,
  input  [63:0] io_ins_407,
  input  [63:0] io_ins_408,
  input  [63:0] io_ins_409,
  input  [63:0] io_ins_410,
  input  [63:0] io_ins_411,
  input  [63:0] io_ins_412,
  input  [63:0] io_ins_413,
  input  [63:0] io_ins_414,
  input  [63:0] io_ins_415,
  input  [63:0] io_ins_416,
  input  [63:0] io_ins_417,
  input  [63:0] io_ins_418,
  input  [63:0] io_ins_419,
  input  [63:0] io_ins_420,
  input  [63:0] io_ins_421,
  input  [63:0] io_ins_422,
  input  [63:0] io_ins_423,
  input  [63:0] io_ins_424,
  input  [63:0] io_ins_425,
  input  [63:0] io_ins_426,
  input  [63:0] io_ins_427,
  input  [63:0] io_ins_428,
  input  [63:0] io_ins_429,
  input  [63:0] io_ins_430,
  input  [63:0] io_ins_431,
  input  [63:0] io_ins_432,
  input  [63:0] io_ins_433,
  input  [63:0] io_ins_434,
  input  [63:0] io_ins_435,
  input  [63:0] io_ins_436,
  input  [63:0] io_ins_437,
  input  [63:0] io_ins_438,
  input  [63:0] io_ins_439,
  input  [63:0] io_ins_440,
  input  [63:0] io_ins_441,
  input  [63:0] io_ins_442,
  input  [63:0] io_ins_443,
  input  [63:0] io_ins_444,
  input  [63:0] io_ins_445,
  input  [63:0] io_ins_446,
  input  [63:0] io_ins_447,
  input  [63:0] io_ins_448,
  input  [63:0] io_ins_449,
  input  [63:0] io_ins_450,
  input  [63:0] io_ins_451,
  input  [63:0] io_ins_452,
  input  [63:0] io_ins_453,
  input  [63:0] io_ins_454,
  input  [63:0] io_ins_455,
  input  [63:0] io_ins_456,
  input  [63:0] io_ins_457,
  input  [63:0] io_ins_458,
  input  [63:0] io_ins_459,
  input  [63:0] io_ins_460,
  input  [63:0] io_ins_461,
  input  [63:0] io_ins_462,
  input  [63:0] io_ins_463,
  input  [63:0] io_ins_464,
  input  [63:0] io_ins_465,
  input  [63:0] io_ins_466,
  input  [63:0] io_ins_467,
  input  [63:0] io_ins_468,
  input  [63:0] io_ins_469,
  input  [63:0] io_ins_470,
  input  [63:0] io_ins_471,
  input  [63:0] io_ins_472,
  input  [63:0] io_ins_473,
  input  [63:0] io_ins_474,
  input  [63:0] io_ins_475,
  input  [63:0] io_ins_476,
  input  [63:0] io_ins_477,
  input  [63:0] io_ins_478,
  input  [63:0] io_ins_479,
  input  [63:0] io_ins_480,
  input  [63:0] io_ins_481,
  input  [63:0] io_ins_482,
  input  [63:0] io_ins_483,
  input  [63:0] io_ins_484,
  input  [63:0] io_ins_485,
  input  [63:0] io_ins_486,
  input  [63:0] io_ins_487,
  input  [63:0] io_ins_488,
  input  [63:0] io_ins_489,
  input  [63:0] io_ins_490,
  input  [63:0] io_ins_491,
  input  [63:0] io_ins_492,
  input  [63:0] io_ins_493,
  input  [63:0] io_ins_494,
  input  [63:0] io_ins_495,
  input  [63:0] io_ins_496,
  input  [63:0] io_ins_497,
  input  [63:0] io_ins_498,
  input  [63:0] io_ins_499,
  input  [63:0] io_ins_500,
  input  [63:0] io_ins_501,
  input  [63:0] io_ins_502,
  input  [63:0] io_ins_503,
  input  [63:0] io_ins_504,
  input  [63:0] io_ins_505,
  input  [8:0]  io_sel,
  output [63:0] io_out
);
  wire [63:0] _GEN_0;
  wire [63:0] _GEN_1;
  wire [63:0] _GEN_2;
  wire [63:0] _GEN_3;
  wire [63:0] _GEN_4;
  wire [63:0] _GEN_5;
  wire [63:0] _GEN_6;
  wire [63:0] _GEN_7;
  wire [63:0] _GEN_8;
  wire [63:0] _GEN_9;
  wire [63:0] _GEN_10;
  wire [63:0] _GEN_11;
  wire [63:0] _GEN_12;
  wire [63:0] _GEN_13;
  wire [63:0] _GEN_14;
  wire [63:0] _GEN_15;
  wire [63:0] _GEN_16;
  wire [63:0] _GEN_17;
  wire [63:0] _GEN_18;
  wire [63:0] _GEN_19;
  wire [63:0] _GEN_20;
  wire [63:0] _GEN_21;
  wire [63:0] _GEN_22;
  wire [63:0] _GEN_23;
  wire [63:0] _GEN_24;
  wire [63:0] _GEN_25;
  wire [63:0] _GEN_26;
  wire [63:0] _GEN_27;
  wire [63:0] _GEN_28;
  wire [63:0] _GEN_29;
  wire [63:0] _GEN_30;
  wire [63:0] _GEN_31;
  wire [63:0] _GEN_32;
  wire [63:0] _GEN_33;
  wire [63:0] _GEN_34;
  wire [63:0] _GEN_35;
  wire [63:0] _GEN_36;
  wire [63:0] _GEN_37;
  wire [63:0] _GEN_38;
  wire [63:0] _GEN_39;
  wire [63:0] _GEN_40;
  wire [63:0] _GEN_41;
  wire [63:0] _GEN_42;
  wire [63:0] _GEN_43;
  wire [63:0] _GEN_44;
  wire [63:0] _GEN_45;
  wire [63:0] _GEN_46;
  wire [63:0] _GEN_47;
  wire [63:0] _GEN_48;
  wire [63:0] _GEN_49;
  wire [63:0] _GEN_50;
  wire [63:0] _GEN_51;
  wire [63:0] _GEN_52;
  wire [63:0] _GEN_53;
  wire [63:0] _GEN_54;
  wire [63:0] _GEN_55;
  wire [63:0] _GEN_56;
  wire [63:0] _GEN_57;
  wire [63:0] _GEN_58;
  wire [63:0] _GEN_59;
  wire [63:0] _GEN_60;
  wire [63:0] _GEN_61;
  wire [63:0] _GEN_62;
  wire [63:0] _GEN_63;
  wire [63:0] _GEN_64;
  wire [63:0] _GEN_65;
  wire [63:0] _GEN_66;
  wire [63:0] _GEN_67;
  wire [63:0] _GEN_68;
  wire [63:0] _GEN_69;
  wire [63:0] _GEN_70;
  wire [63:0] _GEN_71;
  wire [63:0] _GEN_72;
  wire [63:0] _GEN_73;
  wire [63:0] _GEN_74;
  wire [63:0] _GEN_75;
  wire [63:0] _GEN_76;
  wire [63:0] _GEN_77;
  wire [63:0] _GEN_78;
  wire [63:0] _GEN_79;
  wire [63:0] _GEN_80;
  wire [63:0] _GEN_81;
  wire [63:0] _GEN_82;
  wire [63:0] _GEN_83;
  wire [63:0] _GEN_84;
  wire [63:0] _GEN_85;
  wire [63:0] _GEN_86;
  wire [63:0] _GEN_87;
  wire [63:0] _GEN_88;
  wire [63:0] _GEN_89;
  wire [63:0] _GEN_90;
  wire [63:0] _GEN_91;
  wire [63:0] _GEN_92;
  wire [63:0] _GEN_93;
  wire [63:0] _GEN_94;
  wire [63:0] _GEN_95;
  wire [63:0] _GEN_96;
  wire [63:0] _GEN_97;
  wire [63:0] _GEN_98;
  wire [63:0] _GEN_99;
  wire [63:0] _GEN_100;
  wire [63:0] _GEN_101;
  wire [63:0] _GEN_102;
  wire [63:0] _GEN_103;
  wire [63:0] _GEN_104;
  wire [63:0] _GEN_105;
  wire [63:0] _GEN_106;
  wire [63:0] _GEN_107;
  wire [63:0] _GEN_108;
  wire [63:0] _GEN_109;
  wire [63:0] _GEN_110;
  wire [63:0] _GEN_111;
  wire [63:0] _GEN_112;
  wire [63:0] _GEN_113;
  wire [63:0] _GEN_114;
  wire [63:0] _GEN_115;
  wire [63:0] _GEN_116;
  wire [63:0] _GEN_117;
  wire [63:0] _GEN_118;
  wire [63:0] _GEN_119;
  wire [63:0] _GEN_120;
  wire [63:0] _GEN_121;
  wire [63:0] _GEN_122;
  wire [63:0] _GEN_123;
  wire [63:0] _GEN_124;
  wire [63:0] _GEN_125;
  wire [63:0] _GEN_126;
  wire [63:0] _GEN_127;
  wire [63:0] _GEN_128;
  wire [63:0] _GEN_129;
  wire [63:0] _GEN_130;
  wire [63:0] _GEN_131;
  wire [63:0] _GEN_132;
  wire [63:0] _GEN_133;
  wire [63:0] _GEN_134;
  wire [63:0] _GEN_135;
  wire [63:0] _GEN_136;
  wire [63:0] _GEN_137;
  wire [63:0] _GEN_138;
  wire [63:0] _GEN_139;
  wire [63:0] _GEN_140;
  wire [63:0] _GEN_141;
  wire [63:0] _GEN_142;
  wire [63:0] _GEN_143;
  wire [63:0] _GEN_144;
  wire [63:0] _GEN_145;
  wire [63:0] _GEN_146;
  wire [63:0] _GEN_147;
  wire [63:0] _GEN_148;
  wire [63:0] _GEN_149;
  wire [63:0] _GEN_150;
  wire [63:0] _GEN_151;
  wire [63:0] _GEN_152;
  wire [63:0] _GEN_153;
  wire [63:0] _GEN_154;
  wire [63:0] _GEN_155;
  wire [63:0] _GEN_156;
  wire [63:0] _GEN_157;
  wire [63:0] _GEN_158;
  wire [63:0] _GEN_159;
  wire [63:0] _GEN_160;
  wire [63:0] _GEN_161;
  wire [63:0] _GEN_162;
  wire [63:0] _GEN_163;
  wire [63:0] _GEN_164;
  wire [63:0] _GEN_165;
  wire [63:0] _GEN_166;
  wire [63:0] _GEN_167;
  wire [63:0] _GEN_168;
  wire [63:0] _GEN_169;
  wire [63:0] _GEN_170;
  wire [63:0] _GEN_171;
  wire [63:0] _GEN_172;
  wire [63:0] _GEN_173;
  wire [63:0] _GEN_174;
  wire [63:0] _GEN_175;
  wire [63:0] _GEN_176;
  wire [63:0] _GEN_177;
  wire [63:0] _GEN_178;
  wire [63:0] _GEN_179;
  wire [63:0] _GEN_180;
  wire [63:0] _GEN_181;
  wire [63:0] _GEN_182;
  wire [63:0] _GEN_183;
  wire [63:0] _GEN_184;
  wire [63:0] _GEN_185;
  wire [63:0] _GEN_186;
  wire [63:0] _GEN_187;
  wire [63:0] _GEN_188;
  wire [63:0] _GEN_189;
  wire [63:0] _GEN_190;
  wire [63:0] _GEN_191;
  wire [63:0] _GEN_192;
  wire [63:0] _GEN_193;
  wire [63:0] _GEN_194;
  wire [63:0] _GEN_195;
  wire [63:0] _GEN_196;
  wire [63:0] _GEN_197;
  wire [63:0] _GEN_198;
  wire [63:0] _GEN_199;
  wire [63:0] _GEN_200;
  wire [63:0] _GEN_201;
  wire [63:0] _GEN_202;
  wire [63:0] _GEN_203;
  wire [63:0] _GEN_204;
  wire [63:0] _GEN_205;
  wire [63:0] _GEN_206;
  wire [63:0] _GEN_207;
  wire [63:0] _GEN_208;
  wire [63:0] _GEN_209;
  wire [63:0] _GEN_210;
  wire [63:0] _GEN_211;
  wire [63:0] _GEN_212;
  wire [63:0] _GEN_213;
  wire [63:0] _GEN_214;
  wire [63:0] _GEN_215;
  wire [63:0] _GEN_216;
  wire [63:0] _GEN_217;
  wire [63:0] _GEN_218;
  wire [63:0] _GEN_219;
  wire [63:0] _GEN_220;
  wire [63:0] _GEN_221;
  wire [63:0] _GEN_222;
  wire [63:0] _GEN_223;
  wire [63:0] _GEN_224;
  wire [63:0] _GEN_225;
  wire [63:0] _GEN_226;
  wire [63:0] _GEN_227;
  wire [63:0] _GEN_228;
  wire [63:0] _GEN_229;
  wire [63:0] _GEN_230;
  wire [63:0] _GEN_231;
  wire [63:0] _GEN_232;
  wire [63:0] _GEN_233;
  wire [63:0] _GEN_234;
  wire [63:0] _GEN_235;
  wire [63:0] _GEN_236;
  wire [63:0] _GEN_237;
  wire [63:0] _GEN_238;
  wire [63:0] _GEN_239;
  wire [63:0] _GEN_240;
  wire [63:0] _GEN_241;
  wire [63:0] _GEN_242;
  wire [63:0] _GEN_243;
  wire [63:0] _GEN_244;
  wire [63:0] _GEN_245;
  wire [63:0] _GEN_246;
  wire [63:0] _GEN_247;
  wire [63:0] _GEN_248;
  wire [63:0] _GEN_249;
  wire [63:0] _GEN_250;
  wire [63:0] _GEN_251;
  wire [63:0] _GEN_252;
  wire [63:0] _GEN_253;
  wire [63:0] _GEN_254;
  wire [63:0] _GEN_255;
  wire [63:0] _GEN_256;
  wire [63:0] _GEN_257;
  wire [63:0] _GEN_258;
  wire [63:0] _GEN_259;
  wire [63:0] _GEN_260;
  wire [63:0] _GEN_261;
  wire [63:0] _GEN_262;
  wire [63:0] _GEN_263;
  wire [63:0] _GEN_264;
  wire [63:0] _GEN_265;
  wire [63:0] _GEN_266;
  wire [63:0] _GEN_267;
  wire [63:0] _GEN_268;
  wire [63:0] _GEN_269;
  wire [63:0] _GEN_270;
  wire [63:0] _GEN_271;
  wire [63:0] _GEN_272;
  wire [63:0] _GEN_273;
  wire [63:0] _GEN_274;
  wire [63:0] _GEN_275;
  wire [63:0] _GEN_276;
  wire [63:0] _GEN_277;
  wire [63:0] _GEN_278;
  wire [63:0] _GEN_279;
  wire [63:0] _GEN_280;
  wire [63:0] _GEN_281;
  wire [63:0] _GEN_282;
  wire [63:0] _GEN_283;
  wire [63:0] _GEN_284;
  wire [63:0] _GEN_285;
  wire [63:0] _GEN_286;
  wire [63:0] _GEN_287;
  wire [63:0] _GEN_288;
  wire [63:0] _GEN_289;
  wire [63:0] _GEN_290;
  wire [63:0] _GEN_291;
  wire [63:0] _GEN_292;
  wire [63:0] _GEN_293;
  wire [63:0] _GEN_294;
  wire [63:0] _GEN_295;
  wire [63:0] _GEN_296;
  wire [63:0] _GEN_297;
  wire [63:0] _GEN_298;
  wire [63:0] _GEN_299;
  wire [63:0] _GEN_300;
  wire [63:0] _GEN_301;
  wire [63:0] _GEN_302;
  wire [63:0] _GEN_303;
  wire [63:0] _GEN_304;
  wire [63:0] _GEN_305;
  wire [63:0] _GEN_306;
  wire [63:0] _GEN_307;
  wire [63:0] _GEN_308;
  wire [63:0] _GEN_309;
  wire [63:0] _GEN_310;
  wire [63:0] _GEN_311;
  wire [63:0] _GEN_312;
  wire [63:0] _GEN_313;
  wire [63:0] _GEN_314;
  wire [63:0] _GEN_315;
  wire [63:0] _GEN_316;
  wire [63:0] _GEN_317;
  wire [63:0] _GEN_318;
  wire [63:0] _GEN_319;
  wire [63:0] _GEN_320;
  wire [63:0] _GEN_321;
  wire [63:0] _GEN_322;
  wire [63:0] _GEN_323;
  wire [63:0] _GEN_324;
  wire [63:0] _GEN_325;
  wire [63:0] _GEN_326;
  wire [63:0] _GEN_327;
  wire [63:0] _GEN_328;
  wire [63:0] _GEN_329;
  wire [63:0] _GEN_330;
  wire [63:0] _GEN_331;
  wire [63:0] _GEN_332;
  wire [63:0] _GEN_333;
  wire [63:0] _GEN_334;
  wire [63:0] _GEN_335;
  wire [63:0] _GEN_336;
  wire [63:0] _GEN_337;
  wire [63:0] _GEN_338;
  wire [63:0] _GEN_339;
  wire [63:0] _GEN_340;
  wire [63:0] _GEN_341;
  wire [63:0] _GEN_342;
  wire [63:0] _GEN_343;
  wire [63:0] _GEN_344;
  wire [63:0] _GEN_345;
  wire [63:0] _GEN_346;
  wire [63:0] _GEN_347;
  wire [63:0] _GEN_348;
  wire [63:0] _GEN_349;
  wire [63:0] _GEN_350;
  wire [63:0] _GEN_351;
  wire [63:0] _GEN_352;
  wire [63:0] _GEN_353;
  wire [63:0] _GEN_354;
  wire [63:0] _GEN_355;
  wire [63:0] _GEN_356;
  wire [63:0] _GEN_357;
  wire [63:0] _GEN_358;
  wire [63:0] _GEN_359;
  wire [63:0] _GEN_360;
  wire [63:0] _GEN_361;
  wire [63:0] _GEN_362;
  wire [63:0] _GEN_363;
  wire [63:0] _GEN_364;
  wire [63:0] _GEN_365;
  wire [63:0] _GEN_366;
  wire [63:0] _GEN_367;
  wire [63:0] _GEN_368;
  wire [63:0] _GEN_369;
  wire [63:0] _GEN_370;
  wire [63:0] _GEN_371;
  wire [63:0] _GEN_372;
  wire [63:0] _GEN_373;
  wire [63:0] _GEN_374;
  wire [63:0] _GEN_375;
  wire [63:0] _GEN_376;
  wire [63:0] _GEN_377;
  wire [63:0] _GEN_378;
  wire [63:0] _GEN_379;
  wire [63:0] _GEN_380;
  wire [63:0] _GEN_381;
  wire [63:0] _GEN_382;
  wire [63:0] _GEN_383;
  wire [63:0] _GEN_384;
  wire [63:0] _GEN_385;
  wire [63:0] _GEN_386;
  wire [63:0] _GEN_387;
  wire [63:0] _GEN_388;
  wire [63:0] _GEN_389;
  wire [63:0] _GEN_390;
  wire [63:0] _GEN_391;
  wire [63:0] _GEN_392;
  wire [63:0] _GEN_393;
  wire [63:0] _GEN_394;
  wire [63:0] _GEN_395;
  wire [63:0] _GEN_396;
  wire [63:0] _GEN_397;
  wire [63:0] _GEN_398;
  wire [63:0] _GEN_399;
  wire [63:0] _GEN_400;
  wire [63:0] _GEN_401;
  wire [63:0] _GEN_402;
  wire [63:0] _GEN_403;
  wire [63:0] _GEN_404;
  wire [63:0] _GEN_405;
  wire [63:0] _GEN_406;
  wire [63:0] _GEN_407;
  wire [63:0] _GEN_408;
  wire [63:0] _GEN_409;
  wire [63:0] _GEN_410;
  wire [63:0] _GEN_411;
  wire [63:0] _GEN_412;
  wire [63:0] _GEN_413;
  wire [63:0] _GEN_414;
  wire [63:0] _GEN_415;
  wire [63:0] _GEN_416;
  wire [63:0] _GEN_417;
  wire [63:0] _GEN_418;
  wire [63:0] _GEN_419;
  wire [63:0] _GEN_420;
  wire [63:0] _GEN_421;
  wire [63:0] _GEN_422;
  wire [63:0] _GEN_423;
  wire [63:0] _GEN_424;
  wire [63:0] _GEN_425;
  wire [63:0] _GEN_426;
  wire [63:0] _GEN_427;
  wire [63:0] _GEN_428;
  wire [63:0] _GEN_429;
  wire [63:0] _GEN_430;
  wire [63:0] _GEN_431;
  wire [63:0] _GEN_432;
  wire [63:0] _GEN_433;
  wire [63:0] _GEN_434;
  wire [63:0] _GEN_435;
  wire [63:0] _GEN_436;
  wire [63:0] _GEN_437;
  wire [63:0] _GEN_438;
  wire [63:0] _GEN_439;
  wire [63:0] _GEN_440;
  wire [63:0] _GEN_441;
  wire [63:0] _GEN_442;
  wire [63:0] _GEN_443;
  wire [63:0] _GEN_444;
  wire [63:0] _GEN_445;
  wire [63:0] _GEN_446;
  wire [63:0] _GEN_447;
  wire [63:0] _GEN_448;
  wire [63:0] _GEN_449;
  wire [63:0] _GEN_450;
  wire [63:0] _GEN_451;
  wire [63:0] _GEN_452;
  wire [63:0] _GEN_453;
  wire [63:0] _GEN_454;
  wire [63:0] _GEN_455;
  wire [63:0] _GEN_456;
  wire [63:0] _GEN_457;
  wire [63:0] _GEN_458;
  wire [63:0] _GEN_459;
  wire [63:0] _GEN_460;
  wire [63:0] _GEN_461;
  wire [63:0] _GEN_462;
  wire [63:0] _GEN_463;
  wire [63:0] _GEN_464;
  wire [63:0] _GEN_465;
  wire [63:0] _GEN_466;
  wire [63:0] _GEN_467;
  wire [63:0] _GEN_468;
  wire [63:0] _GEN_469;
  wire [63:0] _GEN_470;
  wire [63:0] _GEN_471;
  wire [63:0] _GEN_472;
  wire [63:0] _GEN_473;
  wire [63:0] _GEN_474;
  wire [63:0] _GEN_475;
  wire [63:0] _GEN_476;
  wire [63:0] _GEN_477;
  wire [63:0] _GEN_478;
  wire [63:0] _GEN_479;
  wire [63:0] _GEN_480;
  wire [63:0] _GEN_481;
  wire [63:0] _GEN_482;
  wire [63:0] _GEN_483;
  wire [63:0] _GEN_484;
  wire [63:0] _GEN_485;
  wire [63:0] _GEN_486;
  wire [63:0] _GEN_487;
  wire [63:0] _GEN_488;
  wire [63:0] _GEN_489;
  wire [63:0] _GEN_490;
  wire [63:0] _GEN_491;
  wire [63:0] _GEN_492;
  wire [63:0] _GEN_493;
  wire [63:0] _GEN_494;
  wire [63:0] _GEN_495;
  wire [63:0] _GEN_496;
  wire [63:0] _GEN_497;
  wire [63:0] _GEN_498;
  wire [63:0] _GEN_499;
  wire [63:0] _GEN_500;
  wire [63:0] _GEN_501;
  wire [63:0] _GEN_502;
  wire [63:0] _GEN_503;
  wire [63:0] _GEN_504;
  wire [63:0] _GEN_505;
  assign _GEN_1 = 9'h1 == io_sel ? io_ins_1 : io_ins_0;
  assign _GEN_2 = 9'h2 == io_sel ? io_ins_2 : _GEN_1;
  assign _GEN_3 = 9'h3 == io_sel ? io_ins_3 : _GEN_2;
  assign _GEN_4 = 9'h4 == io_sel ? io_ins_4 : _GEN_3;
  assign _GEN_5 = 9'h5 == io_sel ? io_ins_5 : _GEN_4;
  assign _GEN_6 = 9'h6 == io_sel ? io_ins_6 : _GEN_5;
  assign _GEN_7 = 9'h7 == io_sel ? io_ins_7 : _GEN_6;
  assign _GEN_8 = 9'h8 == io_sel ? io_ins_8 : _GEN_7;
  assign _GEN_9 = 9'h9 == io_sel ? io_ins_9 : _GEN_8;
  assign _GEN_10 = 9'ha == io_sel ? io_ins_10 : _GEN_9;
  assign _GEN_11 = 9'hb == io_sel ? io_ins_11 : _GEN_10;
  assign _GEN_12 = 9'hc == io_sel ? io_ins_12 : _GEN_11;
  assign _GEN_13 = 9'hd == io_sel ? io_ins_13 : _GEN_12;
  assign _GEN_14 = 9'he == io_sel ? io_ins_14 : _GEN_13;
  assign _GEN_15 = 9'hf == io_sel ? io_ins_15 : _GEN_14;
  assign _GEN_16 = 9'h10 == io_sel ? io_ins_16 : _GEN_15;
  assign _GEN_17 = 9'h11 == io_sel ? io_ins_17 : _GEN_16;
  assign _GEN_18 = 9'h12 == io_sel ? io_ins_18 : _GEN_17;
  assign _GEN_19 = 9'h13 == io_sel ? io_ins_19 : _GEN_18;
  assign _GEN_20 = 9'h14 == io_sel ? io_ins_20 : _GEN_19;
  assign _GEN_21 = 9'h15 == io_sel ? io_ins_21 : _GEN_20;
  assign _GEN_22 = 9'h16 == io_sel ? io_ins_22 : _GEN_21;
  assign _GEN_23 = 9'h17 == io_sel ? io_ins_23 : _GEN_22;
  assign _GEN_24 = 9'h18 == io_sel ? io_ins_24 : _GEN_23;
  assign _GEN_25 = 9'h19 == io_sel ? io_ins_25 : _GEN_24;
  assign _GEN_26 = 9'h1a == io_sel ? io_ins_26 : _GEN_25;
  assign _GEN_27 = 9'h1b == io_sel ? io_ins_27 : _GEN_26;
  assign _GEN_28 = 9'h1c == io_sel ? io_ins_28 : _GEN_27;
  assign _GEN_29 = 9'h1d == io_sel ? io_ins_29 : _GEN_28;
  assign _GEN_30 = 9'h1e == io_sel ? io_ins_30 : _GEN_29;
  assign _GEN_31 = 9'h1f == io_sel ? io_ins_31 : _GEN_30;
  assign _GEN_32 = 9'h20 == io_sel ? io_ins_32 : _GEN_31;
  assign _GEN_33 = 9'h21 == io_sel ? io_ins_33 : _GEN_32;
  assign _GEN_34 = 9'h22 == io_sel ? io_ins_34 : _GEN_33;
  assign _GEN_35 = 9'h23 == io_sel ? io_ins_35 : _GEN_34;
  assign _GEN_36 = 9'h24 == io_sel ? io_ins_36 : _GEN_35;
  assign _GEN_37 = 9'h25 == io_sel ? io_ins_37 : _GEN_36;
  assign _GEN_38 = 9'h26 == io_sel ? io_ins_38 : _GEN_37;
  assign _GEN_39 = 9'h27 == io_sel ? io_ins_39 : _GEN_38;
  assign _GEN_40 = 9'h28 == io_sel ? io_ins_40 : _GEN_39;
  assign _GEN_41 = 9'h29 == io_sel ? io_ins_41 : _GEN_40;
  assign _GEN_42 = 9'h2a == io_sel ? io_ins_42 : _GEN_41;
  assign _GEN_43 = 9'h2b == io_sel ? io_ins_43 : _GEN_42;
  assign _GEN_44 = 9'h2c == io_sel ? io_ins_44 : _GEN_43;
  assign _GEN_45 = 9'h2d == io_sel ? io_ins_45 : _GEN_44;
  assign _GEN_46 = 9'h2e == io_sel ? io_ins_46 : _GEN_45;
  assign _GEN_47 = 9'h2f == io_sel ? io_ins_47 : _GEN_46;
  assign _GEN_48 = 9'h30 == io_sel ? io_ins_48 : _GEN_47;
  assign _GEN_49 = 9'h31 == io_sel ? io_ins_49 : _GEN_48;
  assign _GEN_50 = 9'h32 == io_sel ? io_ins_50 : _GEN_49;
  assign _GEN_51 = 9'h33 == io_sel ? io_ins_51 : _GEN_50;
  assign _GEN_52 = 9'h34 == io_sel ? io_ins_52 : _GEN_51;
  assign _GEN_53 = 9'h35 == io_sel ? io_ins_53 : _GEN_52;
  assign _GEN_54 = 9'h36 == io_sel ? io_ins_54 : _GEN_53;
  assign _GEN_55 = 9'h37 == io_sel ? io_ins_55 : _GEN_54;
  assign _GEN_56 = 9'h38 == io_sel ? io_ins_56 : _GEN_55;
  assign _GEN_57 = 9'h39 == io_sel ? io_ins_57 : _GEN_56;
  assign _GEN_58 = 9'h3a == io_sel ? io_ins_58 : _GEN_57;
  assign _GEN_59 = 9'h3b == io_sel ? io_ins_59 : _GEN_58;
  assign _GEN_60 = 9'h3c == io_sel ? io_ins_60 : _GEN_59;
  assign _GEN_61 = 9'h3d == io_sel ? io_ins_61 : _GEN_60;
  assign _GEN_62 = 9'h3e == io_sel ? io_ins_62 : _GEN_61;
  assign _GEN_63 = 9'h3f == io_sel ? io_ins_63 : _GEN_62;
  assign _GEN_64 = 9'h40 == io_sel ? io_ins_64 : _GEN_63;
  assign _GEN_65 = 9'h41 == io_sel ? io_ins_65 : _GEN_64;
  assign _GEN_66 = 9'h42 == io_sel ? io_ins_66 : _GEN_65;
  assign _GEN_67 = 9'h43 == io_sel ? io_ins_67 : _GEN_66;
  assign _GEN_68 = 9'h44 == io_sel ? io_ins_68 : _GEN_67;
  assign _GEN_69 = 9'h45 == io_sel ? io_ins_69 : _GEN_68;
  assign _GEN_70 = 9'h46 == io_sel ? io_ins_70 : _GEN_69;
  assign _GEN_71 = 9'h47 == io_sel ? io_ins_71 : _GEN_70;
  assign _GEN_72 = 9'h48 == io_sel ? io_ins_72 : _GEN_71;
  assign _GEN_73 = 9'h49 == io_sel ? io_ins_73 : _GEN_72;
  assign _GEN_74 = 9'h4a == io_sel ? io_ins_74 : _GEN_73;
  assign _GEN_75 = 9'h4b == io_sel ? io_ins_75 : _GEN_74;
  assign _GEN_76 = 9'h4c == io_sel ? io_ins_76 : _GEN_75;
  assign _GEN_77 = 9'h4d == io_sel ? io_ins_77 : _GEN_76;
  assign _GEN_78 = 9'h4e == io_sel ? io_ins_78 : _GEN_77;
  assign _GEN_79 = 9'h4f == io_sel ? io_ins_79 : _GEN_78;
  assign _GEN_80 = 9'h50 == io_sel ? io_ins_80 : _GEN_79;
  assign _GEN_81 = 9'h51 == io_sel ? io_ins_81 : _GEN_80;
  assign _GEN_82 = 9'h52 == io_sel ? io_ins_82 : _GEN_81;
  assign _GEN_83 = 9'h53 == io_sel ? io_ins_83 : _GEN_82;
  assign _GEN_84 = 9'h54 == io_sel ? io_ins_84 : _GEN_83;
  assign _GEN_85 = 9'h55 == io_sel ? io_ins_85 : _GEN_84;
  assign _GEN_86 = 9'h56 == io_sel ? io_ins_86 : _GEN_85;
  assign _GEN_87 = 9'h57 == io_sel ? io_ins_87 : _GEN_86;
  assign _GEN_88 = 9'h58 == io_sel ? io_ins_88 : _GEN_87;
  assign _GEN_89 = 9'h59 == io_sel ? io_ins_89 : _GEN_88;
  assign _GEN_90 = 9'h5a == io_sel ? io_ins_90 : _GEN_89;
  assign _GEN_91 = 9'h5b == io_sel ? io_ins_91 : _GEN_90;
  assign _GEN_92 = 9'h5c == io_sel ? io_ins_92 : _GEN_91;
  assign _GEN_93 = 9'h5d == io_sel ? io_ins_93 : _GEN_92;
  assign _GEN_94 = 9'h5e == io_sel ? io_ins_94 : _GEN_93;
  assign _GEN_95 = 9'h5f == io_sel ? io_ins_95 : _GEN_94;
  assign _GEN_96 = 9'h60 == io_sel ? io_ins_96 : _GEN_95;
  assign _GEN_97 = 9'h61 == io_sel ? io_ins_97 : _GEN_96;
  assign _GEN_98 = 9'h62 == io_sel ? io_ins_98 : _GEN_97;
  assign _GEN_99 = 9'h63 == io_sel ? io_ins_99 : _GEN_98;
  assign _GEN_100 = 9'h64 == io_sel ? io_ins_100 : _GEN_99;
  assign _GEN_101 = 9'h65 == io_sel ? io_ins_101 : _GEN_100;
  assign _GEN_102 = 9'h66 == io_sel ? io_ins_102 : _GEN_101;
  assign _GEN_103 = 9'h67 == io_sel ? io_ins_103 : _GEN_102;
  assign _GEN_104 = 9'h68 == io_sel ? io_ins_104 : _GEN_103;
  assign _GEN_105 = 9'h69 == io_sel ? io_ins_105 : _GEN_104;
  assign _GEN_106 = 9'h6a == io_sel ? io_ins_106 : _GEN_105;
  assign _GEN_107 = 9'h6b == io_sel ? io_ins_107 : _GEN_106;
  assign _GEN_108 = 9'h6c == io_sel ? io_ins_108 : _GEN_107;
  assign _GEN_109 = 9'h6d == io_sel ? io_ins_109 : _GEN_108;
  assign _GEN_110 = 9'h6e == io_sel ? io_ins_110 : _GEN_109;
  assign _GEN_111 = 9'h6f == io_sel ? io_ins_111 : _GEN_110;
  assign _GEN_112 = 9'h70 == io_sel ? io_ins_112 : _GEN_111;
  assign _GEN_113 = 9'h71 == io_sel ? io_ins_113 : _GEN_112;
  assign _GEN_114 = 9'h72 == io_sel ? io_ins_114 : _GEN_113;
  assign _GEN_115 = 9'h73 == io_sel ? io_ins_115 : _GEN_114;
  assign _GEN_116 = 9'h74 == io_sel ? io_ins_116 : _GEN_115;
  assign _GEN_117 = 9'h75 == io_sel ? io_ins_117 : _GEN_116;
  assign _GEN_118 = 9'h76 == io_sel ? io_ins_118 : _GEN_117;
  assign _GEN_119 = 9'h77 == io_sel ? io_ins_119 : _GEN_118;
  assign _GEN_120 = 9'h78 == io_sel ? io_ins_120 : _GEN_119;
  assign _GEN_121 = 9'h79 == io_sel ? io_ins_121 : _GEN_120;
  assign _GEN_122 = 9'h7a == io_sel ? io_ins_122 : _GEN_121;
  assign _GEN_123 = 9'h7b == io_sel ? io_ins_123 : _GEN_122;
  assign _GEN_124 = 9'h7c == io_sel ? io_ins_124 : _GEN_123;
  assign _GEN_125 = 9'h7d == io_sel ? io_ins_125 : _GEN_124;
  assign _GEN_126 = 9'h7e == io_sel ? io_ins_126 : _GEN_125;
  assign _GEN_127 = 9'h7f == io_sel ? io_ins_127 : _GEN_126;
  assign _GEN_128 = 9'h80 == io_sel ? io_ins_128 : _GEN_127;
  assign _GEN_129 = 9'h81 == io_sel ? io_ins_129 : _GEN_128;
  assign _GEN_130 = 9'h82 == io_sel ? io_ins_130 : _GEN_129;
  assign _GEN_131 = 9'h83 == io_sel ? io_ins_131 : _GEN_130;
  assign _GEN_132 = 9'h84 == io_sel ? io_ins_132 : _GEN_131;
  assign _GEN_133 = 9'h85 == io_sel ? io_ins_133 : _GEN_132;
  assign _GEN_134 = 9'h86 == io_sel ? io_ins_134 : _GEN_133;
  assign _GEN_135 = 9'h87 == io_sel ? io_ins_135 : _GEN_134;
  assign _GEN_136 = 9'h88 == io_sel ? io_ins_136 : _GEN_135;
  assign _GEN_137 = 9'h89 == io_sel ? io_ins_137 : _GEN_136;
  assign _GEN_138 = 9'h8a == io_sel ? io_ins_138 : _GEN_137;
  assign _GEN_139 = 9'h8b == io_sel ? io_ins_139 : _GEN_138;
  assign _GEN_140 = 9'h8c == io_sel ? io_ins_140 : _GEN_139;
  assign _GEN_141 = 9'h8d == io_sel ? io_ins_141 : _GEN_140;
  assign _GEN_142 = 9'h8e == io_sel ? io_ins_142 : _GEN_141;
  assign _GEN_143 = 9'h8f == io_sel ? io_ins_143 : _GEN_142;
  assign _GEN_144 = 9'h90 == io_sel ? io_ins_144 : _GEN_143;
  assign _GEN_145 = 9'h91 == io_sel ? io_ins_145 : _GEN_144;
  assign _GEN_146 = 9'h92 == io_sel ? io_ins_146 : _GEN_145;
  assign _GEN_147 = 9'h93 == io_sel ? io_ins_147 : _GEN_146;
  assign _GEN_148 = 9'h94 == io_sel ? io_ins_148 : _GEN_147;
  assign _GEN_149 = 9'h95 == io_sel ? io_ins_149 : _GEN_148;
  assign _GEN_150 = 9'h96 == io_sel ? io_ins_150 : _GEN_149;
  assign _GEN_151 = 9'h97 == io_sel ? io_ins_151 : _GEN_150;
  assign _GEN_152 = 9'h98 == io_sel ? io_ins_152 : _GEN_151;
  assign _GEN_153 = 9'h99 == io_sel ? io_ins_153 : _GEN_152;
  assign _GEN_154 = 9'h9a == io_sel ? io_ins_154 : _GEN_153;
  assign _GEN_155 = 9'h9b == io_sel ? io_ins_155 : _GEN_154;
  assign _GEN_156 = 9'h9c == io_sel ? io_ins_156 : _GEN_155;
  assign _GEN_157 = 9'h9d == io_sel ? io_ins_157 : _GEN_156;
  assign _GEN_158 = 9'h9e == io_sel ? io_ins_158 : _GEN_157;
  assign _GEN_159 = 9'h9f == io_sel ? io_ins_159 : _GEN_158;
  assign _GEN_160 = 9'ha0 == io_sel ? io_ins_160 : _GEN_159;
  assign _GEN_161 = 9'ha1 == io_sel ? io_ins_161 : _GEN_160;
  assign _GEN_162 = 9'ha2 == io_sel ? io_ins_162 : _GEN_161;
  assign _GEN_163 = 9'ha3 == io_sel ? io_ins_163 : _GEN_162;
  assign _GEN_164 = 9'ha4 == io_sel ? io_ins_164 : _GEN_163;
  assign _GEN_165 = 9'ha5 == io_sel ? io_ins_165 : _GEN_164;
  assign _GEN_166 = 9'ha6 == io_sel ? io_ins_166 : _GEN_165;
  assign _GEN_167 = 9'ha7 == io_sel ? io_ins_167 : _GEN_166;
  assign _GEN_168 = 9'ha8 == io_sel ? io_ins_168 : _GEN_167;
  assign _GEN_169 = 9'ha9 == io_sel ? io_ins_169 : _GEN_168;
  assign _GEN_170 = 9'haa == io_sel ? io_ins_170 : _GEN_169;
  assign _GEN_171 = 9'hab == io_sel ? io_ins_171 : _GEN_170;
  assign _GEN_172 = 9'hac == io_sel ? io_ins_172 : _GEN_171;
  assign _GEN_173 = 9'had == io_sel ? io_ins_173 : _GEN_172;
  assign _GEN_174 = 9'hae == io_sel ? io_ins_174 : _GEN_173;
  assign _GEN_175 = 9'haf == io_sel ? io_ins_175 : _GEN_174;
  assign _GEN_176 = 9'hb0 == io_sel ? io_ins_176 : _GEN_175;
  assign _GEN_177 = 9'hb1 == io_sel ? io_ins_177 : _GEN_176;
  assign _GEN_178 = 9'hb2 == io_sel ? io_ins_178 : _GEN_177;
  assign _GEN_179 = 9'hb3 == io_sel ? io_ins_179 : _GEN_178;
  assign _GEN_180 = 9'hb4 == io_sel ? io_ins_180 : _GEN_179;
  assign _GEN_181 = 9'hb5 == io_sel ? io_ins_181 : _GEN_180;
  assign _GEN_182 = 9'hb6 == io_sel ? io_ins_182 : _GEN_181;
  assign _GEN_183 = 9'hb7 == io_sel ? io_ins_183 : _GEN_182;
  assign _GEN_184 = 9'hb8 == io_sel ? io_ins_184 : _GEN_183;
  assign _GEN_185 = 9'hb9 == io_sel ? io_ins_185 : _GEN_184;
  assign _GEN_186 = 9'hba == io_sel ? io_ins_186 : _GEN_185;
  assign _GEN_187 = 9'hbb == io_sel ? io_ins_187 : _GEN_186;
  assign _GEN_188 = 9'hbc == io_sel ? io_ins_188 : _GEN_187;
  assign _GEN_189 = 9'hbd == io_sel ? io_ins_189 : _GEN_188;
  assign _GEN_190 = 9'hbe == io_sel ? io_ins_190 : _GEN_189;
  assign _GEN_191 = 9'hbf == io_sel ? io_ins_191 : _GEN_190;
  assign _GEN_192 = 9'hc0 == io_sel ? io_ins_192 : _GEN_191;
  assign _GEN_193 = 9'hc1 == io_sel ? io_ins_193 : _GEN_192;
  assign _GEN_194 = 9'hc2 == io_sel ? io_ins_194 : _GEN_193;
  assign _GEN_195 = 9'hc3 == io_sel ? io_ins_195 : _GEN_194;
  assign _GEN_196 = 9'hc4 == io_sel ? io_ins_196 : _GEN_195;
  assign _GEN_197 = 9'hc5 == io_sel ? io_ins_197 : _GEN_196;
  assign _GEN_198 = 9'hc6 == io_sel ? io_ins_198 : _GEN_197;
  assign _GEN_199 = 9'hc7 == io_sel ? io_ins_199 : _GEN_198;
  assign _GEN_200 = 9'hc8 == io_sel ? io_ins_200 : _GEN_199;
  assign _GEN_201 = 9'hc9 == io_sel ? io_ins_201 : _GEN_200;
  assign _GEN_202 = 9'hca == io_sel ? io_ins_202 : _GEN_201;
  assign _GEN_203 = 9'hcb == io_sel ? io_ins_203 : _GEN_202;
  assign _GEN_204 = 9'hcc == io_sel ? io_ins_204 : _GEN_203;
  assign _GEN_205 = 9'hcd == io_sel ? io_ins_205 : _GEN_204;
  assign _GEN_206 = 9'hce == io_sel ? io_ins_206 : _GEN_205;
  assign _GEN_207 = 9'hcf == io_sel ? io_ins_207 : _GEN_206;
  assign _GEN_208 = 9'hd0 == io_sel ? io_ins_208 : _GEN_207;
  assign _GEN_209 = 9'hd1 == io_sel ? io_ins_209 : _GEN_208;
  assign _GEN_210 = 9'hd2 == io_sel ? io_ins_210 : _GEN_209;
  assign _GEN_211 = 9'hd3 == io_sel ? io_ins_211 : _GEN_210;
  assign _GEN_212 = 9'hd4 == io_sel ? io_ins_212 : _GEN_211;
  assign _GEN_213 = 9'hd5 == io_sel ? io_ins_213 : _GEN_212;
  assign _GEN_214 = 9'hd6 == io_sel ? io_ins_214 : _GEN_213;
  assign _GEN_215 = 9'hd7 == io_sel ? io_ins_215 : _GEN_214;
  assign _GEN_216 = 9'hd8 == io_sel ? io_ins_216 : _GEN_215;
  assign _GEN_217 = 9'hd9 == io_sel ? io_ins_217 : _GEN_216;
  assign _GEN_218 = 9'hda == io_sel ? io_ins_218 : _GEN_217;
  assign _GEN_219 = 9'hdb == io_sel ? io_ins_219 : _GEN_218;
  assign _GEN_220 = 9'hdc == io_sel ? io_ins_220 : _GEN_219;
  assign _GEN_221 = 9'hdd == io_sel ? io_ins_221 : _GEN_220;
  assign _GEN_222 = 9'hde == io_sel ? io_ins_222 : _GEN_221;
  assign _GEN_223 = 9'hdf == io_sel ? io_ins_223 : _GEN_222;
  assign _GEN_224 = 9'he0 == io_sel ? io_ins_224 : _GEN_223;
  assign _GEN_225 = 9'he1 == io_sel ? io_ins_225 : _GEN_224;
  assign _GEN_226 = 9'he2 == io_sel ? io_ins_226 : _GEN_225;
  assign _GEN_227 = 9'he3 == io_sel ? io_ins_227 : _GEN_226;
  assign _GEN_228 = 9'he4 == io_sel ? io_ins_228 : _GEN_227;
  assign _GEN_229 = 9'he5 == io_sel ? io_ins_229 : _GEN_228;
  assign _GEN_230 = 9'he6 == io_sel ? io_ins_230 : _GEN_229;
  assign _GEN_231 = 9'he7 == io_sel ? io_ins_231 : _GEN_230;
  assign _GEN_232 = 9'he8 == io_sel ? io_ins_232 : _GEN_231;
  assign _GEN_233 = 9'he9 == io_sel ? io_ins_233 : _GEN_232;
  assign _GEN_234 = 9'hea == io_sel ? io_ins_234 : _GEN_233;
  assign _GEN_235 = 9'heb == io_sel ? io_ins_235 : _GEN_234;
  assign _GEN_236 = 9'hec == io_sel ? io_ins_236 : _GEN_235;
  assign _GEN_237 = 9'hed == io_sel ? io_ins_237 : _GEN_236;
  assign _GEN_238 = 9'hee == io_sel ? io_ins_238 : _GEN_237;
  assign _GEN_239 = 9'hef == io_sel ? io_ins_239 : _GEN_238;
  assign _GEN_240 = 9'hf0 == io_sel ? io_ins_240 : _GEN_239;
  assign _GEN_241 = 9'hf1 == io_sel ? io_ins_241 : _GEN_240;
  assign _GEN_242 = 9'hf2 == io_sel ? io_ins_242 : _GEN_241;
  assign _GEN_243 = 9'hf3 == io_sel ? io_ins_243 : _GEN_242;
  assign _GEN_244 = 9'hf4 == io_sel ? io_ins_244 : _GEN_243;
  assign _GEN_245 = 9'hf5 == io_sel ? io_ins_245 : _GEN_244;
  assign _GEN_246 = 9'hf6 == io_sel ? io_ins_246 : _GEN_245;
  assign _GEN_247 = 9'hf7 == io_sel ? io_ins_247 : _GEN_246;
  assign _GEN_248 = 9'hf8 == io_sel ? io_ins_248 : _GEN_247;
  assign _GEN_249 = 9'hf9 == io_sel ? io_ins_249 : _GEN_248;
  assign _GEN_250 = 9'hfa == io_sel ? io_ins_250 : _GEN_249;
  assign _GEN_251 = 9'hfb == io_sel ? io_ins_251 : _GEN_250;
  assign _GEN_252 = 9'hfc == io_sel ? io_ins_252 : _GEN_251;
  assign _GEN_253 = 9'hfd == io_sel ? io_ins_253 : _GEN_252;
  assign _GEN_254 = 9'hfe == io_sel ? io_ins_254 : _GEN_253;
  assign _GEN_255 = 9'hff == io_sel ? io_ins_255 : _GEN_254;
  assign _GEN_256 = 9'h100 == io_sel ? io_ins_256 : _GEN_255;
  assign _GEN_257 = 9'h101 == io_sel ? io_ins_257 : _GEN_256;
  assign _GEN_258 = 9'h102 == io_sel ? io_ins_258 : _GEN_257;
  assign _GEN_259 = 9'h103 == io_sel ? io_ins_259 : _GEN_258;
  assign _GEN_260 = 9'h104 == io_sel ? io_ins_260 : _GEN_259;
  assign _GEN_261 = 9'h105 == io_sel ? io_ins_261 : _GEN_260;
  assign _GEN_262 = 9'h106 == io_sel ? io_ins_262 : _GEN_261;
  assign _GEN_263 = 9'h107 == io_sel ? io_ins_263 : _GEN_262;
  assign _GEN_264 = 9'h108 == io_sel ? io_ins_264 : _GEN_263;
  assign _GEN_265 = 9'h109 == io_sel ? io_ins_265 : _GEN_264;
  assign _GEN_266 = 9'h10a == io_sel ? io_ins_266 : _GEN_265;
  assign _GEN_267 = 9'h10b == io_sel ? io_ins_267 : _GEN_266;
  assign _GEN_268 = 9'h10c == io_sel ? io_ins_268 : _GEN_267;
  assign _GEN_269 = 9'h10d == io_sel ? io_ins_269 : _GEN_268;
  assign _GEN_270 = 9'h10e == io_sel ? io_ins_270 : _GEN_269;
  assign _GEN_271 = 9'h10f == io_sel ? io_ins_271 : _GEN_270;
  assign _GEN_272 = 9'h110 == io_sel ? io_ins_272 : _GEN_271;
  assign _GEN_273 = 9'h111 == io_sel ? io_ins_273 : _GEN_272;
  assign _GEN_274 = 9'h112 == io_sel ? io_ins_274 : _GEN_273;
  assign _GEN_275 = 9'h113 == io_sel ? io_ins_275 : _GEN_274;
  assign _GEN_276 = 9'h114 == io_sel ? io_ins_276 : _GEN_275;
  assign _GEN_277 = 9'h115 == io_sel ? io_ins_277 : _GEN_276;
  assign _GEN_278 = 9'h116 == io_sel ? io_ins_278 : _GEN_277;
  assign _GEN_279 = 9'h117 == io_sel ? io_ins_279 : _GEN_278;
  assign _GEN_280 = 9'h118 == io_sel ? io_ins_280 : _GEN_279;
  assign _GEN_281 = 9'h119 == io_sel ? io_ins_281 : _GEN_280;
  assign _GEN_282 = 9'h11a == io_sel ? io_ins_282 : _GEN_281;
  assign _GEN_283 = 9'h11b == io_sel ? io_ins_283 : _GEN_282;
  assign _GEN_284 = 9'h11c == io_sel ? io_ins_284 : _GEN_283;
  assign _GEN_285 = 9'h11d == io_sel ? io_ins_285 : _GEN_284;
  assign _GEN_286 = 9'h11e == io_sel ? io_ins_286 : _GEN_285;
  assign _GEN_287 = 9'h11f == io_sel ? io_ins_287 : _GEN_286;
  assign _GEN_288 = 9'h120 == io_sel ? io_ins_288 : _GEN_287;
  assign _GEN_289 = 9'h121 == io_sel ? io_ins_289 : _GEN_288;
  assign _GEN_290 = 9'h122 == io_sel ? io_ins_290 : _GEN_289;
  assign _GEN_291 = 9'h123 == io_sel ? io_ins_291 : _GEN_290;
  assign _GEN_292 = 9'h124 == io_sel ? io_ins_292 : _GEN_291;
  assign _GEN_293 = 9'h125 == io_sel ? io_ins_293 : _GEN_292;
  assign _GEN_294 = 9'h126 == io_sel ? io_ins_294 : _GEN_293;
  assign _GEN_295 = 9'h127 == io_sel ? io_ins_295 : _GEN_294;
  assign _GEN_296 = 9'h128 == io_sel ? io_ins_296 : _GEN_295;
  assign _GEN_297 = 9'h129 == io_sel ? io_ins_297 : _GEN_296;
  assign _GEN_298 = 9'h12a == io_sel ? io_ins_298 : _GEN_297;
  assign _GEN_299 = 9'h12b == io_sel ? io_ins_299 : _GEN_298;
  assign _GEN_300 = 9'h12c == io_sel ? io_ins_300 : _GEN_299;
  assign _GEN_301 = 9'h12d == io_sel ? io_ins_301 : _GEN_300;
  assign _GEN_302 = 9'h12e == io_sel ? io_ins_302 : _GEN_301;
  assign _GEN_303 = 9'h12f == io_sel ? io_ins_303 : _GEN_302;
  assign _GEN_304 = 9'h130 == io_sel ? io_ins_304 : _GEN_303;
  assign _GEN_305 = 9'h131 == io_sel ? io_ins_305 : _GEN_304;
  assign _GEN_306 = 9'h132 == io_sel ? io_ins_306 : _GEN_305;
  assign _GEN_307 = 9'h133 == io_sel ? io_ins_307 : _GEN_306;
  assign _GEN_308 = 9'h134 == io_sel ? io_ins_308 : _GEN_307;
  assign _GEN_309 = 9'h135 == io_sel ? io_ins_309 : _GEN_308;
  assign _GEN_310 = 9'h136 == io_sel ? io_ins_310 : _GEN_309;
  assign _GEN_311 = 9'h137 == io_sel ? io_ins_311 : _GEN_310;
  assign _GEN_312 = 9'h138 == io_sel ? io_ins_312 : _GEN_311;
  assign _GEN_313 = 9'h139 == io_sel ? io_ins_313 : _GEN_312;
  assign _GEN_314 = 9'h13a == io_sel ? io_ins_314 : _GEN_313;
  assign _GEN_315 = 9'h13b == io_sel ? io_ins_315 : _GEN_314;
  assign _GEN_316 = 9'h13c == io_sel ? io_ins_316 : _GEN_315;
  assign _GEN_317 = 9'h13d == io_sel ? io_ins_317 : _GEN_316;
  assign _GEN_318 = 9'h13e == io_sel ? io_ins_318 : _GEN_317;
  assign _GEN_319 = 9'h13f == io_sel ? io_ins_319 : _GEN_318;
  assign _GEN_320 = 9'h140 == io_sel ? io_ins_320 : _GEN_319;
  assign _GEN_321 = 9'h141 == io_sel ? io_ins_321 : _GEN_320;
  assign _GEN_322 = 9'h142 == io_sel ? io_ins_322 : _GEN_321;
  assign _GEN_323 = 9'h143 == io_sel ? io_ins_323 : _GEN_322;
  assign _GEN_324 = 9'h144 == io_sel ? io_ins_324 : _GEN_323;
  assign _GEN_325 = 9'h145 == io_sel ? io_ins_325 : _GEN_324;
  assign _GEN_326 = 9'h146 == io_sel ? io_ins_326 : _GEN_325;
  assign _GEN_327 = 9'h147 == io_sel ? io_ins_327 : _GEN_326;
  assign _GEN_328 = 9'h148 == io_sel ? io_ins_328 : _GEN_327;
  assign _GEN_329 = 9'h149 == io_sel ? io_ins_329 : _GEN_328;
  assign _GEN_330 = 9'h14a == io_sel ? io_ins_330 : _GEN_329;
  assign _GEN_331 = 9'h14b == io_sel ? io_ins_331 : _GEN_330;
  assign _GEN_332 = 9'h14c == io_sel ? io_ins_332 : _GEN_331;
  assign _GEN_333 = 9'h14d == io_sel ? io_ins_333 : _GEN_332;
  assign _GEN_334 = 9'h14e == io_sel ? io_ins_334 : _GEN_333;
  assign _GEN_335 = 9'h14f == io_sel ? io_ins_335 : _GEN_334;
  assign _GEN_336 = 9'h150 == io_sel ? io_ins_336 : _GEN_335;
  assign _GEN_337 = 9'h151 == io_sel ? io_ins_337 : _GEN_336;
  assign _GEN_338 = 9'h152 == io_sel ? io_ins_338 : _GEN_337;
  assign _GEN_339 = 9'h153 == io_sel ? io_ins_339 : _GEN_338;
  assign _GEN_340 = 9'h154 == io_sel ? io_ins_340 : _GEN_339;
  assign _GEN_341 = 9'h155 == io_sel ? io_ins_341 : _GEN_340;
  assign _GEN_342 = 9'h156 == io_sel ? io_ins_342 : _GEN_341;
  assign _GEN_343 = 9'h157 == io_sel ? io_ins_343 : _GEN_342;
  assign _GEN_344 = 9'h158 == io_sel ? io_ins_344 : _GEN_343;
  assign _GEN_345 = 9'h159 == io_sel ? io_ins_345 : _GEN_344;
  assign _GEN_346 = 9'h15a == io_sel ? io_ins_346 : _GEN_345;
  assign _GEN_347 = 9'h15b == io_sel ? io_ins_347 : _GEN_346;
  assign _GEN_348 = 9'h15c == io_sel ? io_ins_348 : _GEN_347;
  assign _GEN_349 = 9'h15d == io_sel ? io_ins_349 : _GEN_348;
  assign _GEN_350 = 9'h15e == io_sel ? io_ins_350 : _GEN_349;
  assign _GEN_351 = 9'h15f == io_sel ? io_ins_351 : _GEN_350;
  assign _GEN_352 = 9'h160 == io_sel ? io_ins_352 : _GEN_351;
  assign _GEN_353 = 9'h161 == io_sel ? io_ins_353 : _GEN_352;
  assign _GEN_354 = 9'h162 == io_sel ? io_ins_354 : _GEN_353;
  assign _GEN_355 = 9'h163 == io_sel ? io_ins_355 : _GEN_354;
  assign _GEN_356 = 9'h164 == io_sel ? io_ins_356 : _GEN_355;
  assign _GEN_357 = 9'h165 == io_sel ? io_ins_357 : _GEN_356;
  assign _GEN_358 = 9'h166 == io_sel ? io_ins_358 : _GEN_357;
  assign _GEN_359 = 9'h167 == io_sel ? io_ins_359 : _GEN_358;
  assign _GEN_360 = 9'h168 == io_sel ? io_ins_360 : _GEN_359;
  assign _GEN_361 = 9'h169 == io_sel ? io_ins_361 : _GEN_360;
  assign _GEN_362 = 9'h16a == io_sel ? io_ins_362 : _GEN_361;
  assign _GEN_363 = 9'h16b == io_sel ? io_ins_363 : _GEN_362;
  assign _GEN_364 = 9'h16c == io_sel ? io_ins_364 : _GEN_363;
  assign _GEN_365 = 9'h16d == io_sel ? io_ins_365 : _GEN_364;
  assign _GEN_366 = 9'h16e == io_sel ? io_ins_366 : _GEN_365;
  assign _GEN_367 = 9'h16f == io_sel ? io_ins_367 : _GEN_366;
  assign _GEN_368 = 9'h170 == io_sel ? io_ins_368 : _GEN_367;
  assign _GEN_369 = 9'h171 == io_sel ? io_ins_369 : _GEN_368;
  assign _GEN_370 = 9'h172 == io_sel ? io_ins_370 : _GEN_369;
  assign _GEN_371 = 9'h173 == io_sel ? io_ins_371 : _GEN_370;
  assign _GEN_372 = 9'h174 == io_sel ? io_ins_372 : _GEN_371;
  assign _GEN_373 = 9'h175 == io_sel ? io_ins_373 : _GEN_372;
  assign _GEN_374 = 9'h176 == io_sel ? io_ins_374 : _GEN_373;
  assign _GEN_375 = 9'h177 == io_sel ? io_ins_375 : _GEN_374;
  assign _GEN_376 = 9'h178 == io_sel ? io_ins_376 : _GEN_375;
  assign _GEN_377 = 9'h179 == io_sel ? io_ins_377 : _GEN_376;
  assign _GEN_378 = 9'h17a == io_sel ? io_ins_378 : _GEN_377;
  assign _GEN_379 = 9'h17b == io_sel ? io_ins_379 : _GEN_378;
  assign _GEN_380 = 9'h17c == io_sel ? io_ins_380 : _GEN_379;
  assign _GEN_381 = 9'h17d == io_sel ? io_ins_381 : _GEN_380;
  assign _GEN_382 = 9'h17e == io_sel ? io_ins_382 : _GEN_381;
  assign _GEN_383 = 9'h17f == io_sel ? io_ins_383 : _GEN_382;
  assign _GEN_384 = 9'h180 == io_sel ? io_ins_384 : _GEN_383;
  assign _GEN_385 = 9'h181 == io_sel ? io_ins_385 : _GEN_384;
  assign _GEN_386 = 9'h182 == io_sel ? io_ins_386 : _GEN_385;
  assign _GEN_387 = 9'h183 == io_sel ? io_ins_387 : _GEN_386;
  assign _GEN_388 = 9'h184 == io_sel ? io_ins_388 : _GEN_387;
  assign _GEN_389 = 9'h185 == io_sel ? io_ins_389 : _GEN_388;
  assign _GEN_390 = 9'h186 == io_sel ? io_ins_390 : _GEN_389;
  assign _GEN_391 = 9'h187 == io_sel ? io_ins_391 : _GEN_390;
  assign _GEN_392 = 9'h188 == io_sel ? io_ins_392 : _GEN_391;
  assign _GEN_393 = 9'h189 == io_sel ? io_ins_393 : _GEN_392;
  assign _GEN_394 = 9'h18a == io_sel ? io_ins_394 : _GEN_393;
  assign _GEN_395 = 9'h18b == io_sel ? io_ins_395 : _GEN_394;
  assign _GEN_396 = 9'h18c == io_sel ? io_ins_396 : _GEN_395;
  assign _GEN_397 = 9'h18d == io_sel ? io_ins_397 : _GEN_396;
  assign _GEN_398 = 9'h18e == io_sel ? io_ins_398 : _GEN_397;
  assign _GEN_399 = 9'h18f == io_sel ? io_ins_399 : _GEN_398;
  assign _GEN_400 = 9'h190 == io_sel ? io_ins_400 : _GEN_399;
  assign _GEN_401 = 9'h191 == io_sel ? io_ins_401 : _GEN_400;
  assign _GEN_402 = 9'h192 == io_sel ? io_ins_402 : _GEN_401;
  assign _GEN_403 = 9'h193 == io_sel ? io_ins_403 : _GEN_402;
  assign _GEN_404 = 9'h194 == io_sel ? io_ins_404 : _GEN_403;
  assign _GEN_405 = 9'h195 == io_sel ? io_ins_405 : _GEN_404;
  assign _GEN_406 = 9'h196 == io_sel ? io_ins_406 : _GEN_405;
  assign _GEN_407 = 9'h197 == io_sel ? io_ins_407 : _GEN_406;
  assign _GEN_408 = 9'h198 == io_sel ? io_ins_408 : _GEN_407;
  assign _GEN_409 = 9'h199 == io_sel ? io_ins_409 : _GEN_408;
  assign _GEN_410 = 9'h19a == io_sel ? io_ins_410 : _GEN_409;
  assign _GEN_411 = 9'h19b == io_sel ? io_ins_411 : _GEN_410;
  assign _GEN_412 = 9'h19c == io_sel ? io_ins_412 : _GEN_411;
  assign _GEN_413 = 9'h19d == io_sel ? io_ins_413 : _GEN_412;
  assign _GEN_414 = 9'h19e == io_sel ? io_ins_414 : _GEN_413;
  assign _GEN_415 = 9'h19f == io_sel ? io_ins_415 : _GEN_414;
  assign _GEN_416 = 9'h1a0 == io_sel ? io_ins_416 : _GEN_415;
  assign _GEN_417 = 9'h1a1 == io_sel ? io_ins_417 : _GEN_416;
  assign _GEN_418 = 9'h1a2 == io_sel ? io_ins_418 : _GEN_417;
  assign _GEN_419 = 9'h1a3 == io_sel ? io_ins_419 : _GEN_418;
  assign _GEN_420 = 9'h1a4 == io_sel ? io_ins_420 : _GEN_419;
  assign _GEN_421 = 9'h1a5 == io_sel ? io_ins_421 : _GEN_420;
  assign _GEN_422 = 9'h1a6 == io_sel ? io_ins_422 : _GEN_421;
  assign _GEN_423 = 9'h1a7 == io_sel ? io_ins_423 : _GEN_422;
  assign _GEN_424 = 9'h1a8 == io_sel ? io_ins_424 : _GEN_423;
  assign _GEN_425 = 9'h1a9 == io_sel ? io_ins_425 : _GEN_424;
  assign _GEN_426 = 9'h1aa == io_sel ? io_ins_426 : _GEN_425;
  assign _GEN_427 = 9'h1ab == io_sel ? io_ins_427 : _GEN_426;
  assign _GEN_428 = 9'h1ac == io_sel ? io_ins_428 : _GEN_427;
  assign _GEN_429 = 9'h1ad == io_sel ? io_ins_429 : _GEN_428;
  assign _GEN_430 = 9'h1ae == io_sel ? io_ins_430 : _GEN_429;
  assign _GEN_431 = 9'h1af == io_sel ? io_ins_431 : _GEN_430;
  assign _GEN_432 = 9'h1b0 == io_sel ? io_ins_432 : _GEN_431;
  assign _GEN_433 = 9'h1b1 == io_sel ? io_ins_433 : _GEN_432;
  assign _GEN_434 = 9'h1b2 == io_sel ? io_ins_434 : _GEN_433;
  assign _GEN_435 = 9'h1b3 == io_sel ? io_ins_435 : _GEN_434;
  assign _GEN_436 = 9'h1b4 == io_sel ? io_ins_436 : _GEN_435;
  assign _GEN_437 = 9'h1b5 == io_sel ? io_ins_437 : _GEN_436;
  assign _GEN_438 = 9'h1b6 == io_sel ? io_ins_438 : _GEN_437;
  assign _GEN_439 = 9'h1b7 == io_sel ? io_ins_439 : _GEN_438;
  assign _GEN_440 = 9'h1b8 == io_sel ? io_ins_440 : _GEN_439;
  assign _GEN_441 = 9'h1b9 == io_sel ? io_ins_441 : _GEN_440;
  assign _GEN_442 = 9'h1ba == io_sel ? io_ins_442 : _GEN_441;
  assign _GEN_443 = 9'h1bb == io_sel ? io_ins_443 : _GEN_442;
  assign _GEN_444 = 9'h1bc == io_sel ? io_ins_444 : _GEN_443;
  assign _GEN_445 = 9'h1bd == io_sel ? io_ins_445 : _GEN_444;
  assign _GEN_446 = 9'h1be == io_sel ? io_ins_446 : _GEN_445;
  assign _GEN_447 = 9'h1bf == io_sel ? io_ins_447 : _GEN_446;
  assign _GEN_448 = 9'h1c0 == io_sel ? io_ins_448 : _GEN_447;
  assign _GEN_449 = 9'h1c1 == io_sel ? io_ins_449 : _GEN_448;
  assign _GEN_450 = 9'h1c2 == io_sel ? io_ins_450 : _GEN_449;
  assign _GEN_451 = 9'h1c3 == io_sel ? io_ins_451 : _GEN_450;
  assign _GEN_452 = 9'h1c4 == io_sel ? io_ins_452 : _GEN_451;
  assign _GEN_453 = 9'h1c5 == io_sel ? io_ins_453 : _GEN_452;
  assign _GEN_454 = 9'h1c6 == io_sel ? io_ins_454 : _GEN_453;
  assign _GEN_455 = 9'h1c7 == io_sel ? io_ins_455 : _GEN_454;
  assign _GEN_456 = 9'h1c8 == io_sel ? io_ins_456 : _GEN_455;
  assign _GEN_457 = 9'h1c9 == io_sel ? io_ins_457 : _GEN_456;
  assign _GEN_458 = 9'h1ca == io_sel ? io_ins_458 : _GEN_457;
  assign _GEN_459 = 9'h1cb == io_sel ? io_ins_459 : _GEN_458;
  assign _GEN_460 = 9'h1cc == io_sel ? io_ins_460 : _GEN_459;
  assign _GEN_461 = 9'h1cd == io_sel ? io_ins_461 : _GEN_460;
  assign _GEN_462 = 9'h1ce == io_sel ? io_ins_462 : _GEN_461;
  assign _GEN_463 = 9'h1cf == io_sel ? io_ins_463 : _GEN_462;
  assign _GEN_464 = 9'h1d0 == io_sel ? io_ins_464 : _GEN_463;
  assign _GEN_465 = 9'h1d1 == io_sel ? io_ins_465 : _GEN_464;
  assign _GEN_466 = 9'h1d2 == io_sel ? io_ins_466 : _GEN_465;
  assign _GEN_467 = 9'h1d3 == io_sel ? io_ins_467 : _GEN_466;
  assign _GEN_468 = 9'h1d4 == io_sel ? io_ins_468 : _GEN_467;
  assign _GEN_469 = 9'h1d5 == io_sel ? io_ins_469 : _GEN_468;
  assign _GEN_470 = 9'h1d6 == io_sel ? io_ins_470 : _GEN_469;
  assign _GEN_471 = 9'h1d7 == io_sel ? io_ins_471 : _GEN_470;
  assign _GEN_472 = 9'h1d8 == io_sel ? io_ins_472 : _GEN_471;
  assign _GEN_473 = 9'h1d9 == io_sel ? io_ins_473 : _GEN_472;
  assign _GEN_474 = 9'h1da == io_sel ? io_ins_474 : _GEN_473;
  assign _GEN_475 = 9'h1db == io_sel ? io_ins_475 : _GEN_474;
  assign _GEN_476 = 9'h1dc == io_sel ? io_ins_476 : _GEN_475;
  assign _GEN_477 = 9'h1dd == io_sel ? io_ins_477 : _GEN_476;
  assign _GEN_478 = 9'h1de == io_sel ? io_ins_478 : _GEN_477;
  assign _GEN_479 = 9'h1df == io_sel ? io_ins_479 : _GEN_478;
  assign _GEN_480 = 9'h1e0 == io_sel ? io_ins_480 : _GEN_479;
  assign _GEN_481 = 9'h1e1 == io_sel ? io_ins_481 : _GEN_480;
  assign _GEN_482 = 9'h1e2 == io_sel ? io_ins_482 : _GEN_481;
  assign _GEN_483 = 9'h1e3 == io_sel ? io_ins_483 : _GEN_482;
  assign _GEN_484 = 9'h1e4 == io_sel ? io_ins_484 : _GEN_483;
  assign _GEN_485 = 9'h1e5 == io_sel ? io_ins_485 : _GEN_484;
  assign _GEN_486 = 9'h1e6 == io_sel ? io_ins_486 : _GEN_485;
  assign _GEN_487 = 9'h1e7 == io_sel ? io_ins_487 : _GEN_486;
  assign _GEN_488 = 9'h1e8 == io_sel ? io_ins_488 : _GEN_487;
  assign _GEN_489 = 9'h1e9 == io_sel ? io_ins_489 : _GEN_488;
  assign _GEN_490 = 9'h1ea == io_sel ? io_ins_490 : _GEN_489;
  assign _GEN_491 = 9'h1eb == io_sel ? io_ins_491 : _GEN_490;
  assign _GEN_492 = 9'h1ec == io_sel ? io_ins_492 : _GEN_491;
  assign _GEN_493 = 9'h1ed == io_sel ? io_ins_493 : _GEN_492;
  assign _GEN_494 = 9'h1ee == io_sel ? io_ins_494 : _GEN_493;
  assign _GEN_495 = 9'h1ef == io_sel ? io_ins_495 : _GEN_494;
  assign _GEN_496 = 9'h1f0 == io_sel ? io_ins_496 : _GEN_495;
  assign _GEN_497 = 9'h1f1 == io_sel ? io_ins_497 : _GEN_496;
  assign _GEN_498 = 9'h1f2 == io_sel ? io_ins_498 : _GEN_497;
  assign _GEN_499 = 9'h1f3 == io_sel ? io_ins_499 : _GEN_498;
  assign _GEN_500 = 9'h1f4 == io_sel ? io_ins_500 : _GEN_499;
  assign _GEN_501 = 9'h1f5 == io_sel ? io_ins_501 : _GEN_500;
  assign _GEN_502 = 9'h1f6 == io_sel ? io_ins_502 : _GEN_501;
  assign _GEN_503 = 9'h1f7 == io_sel ? io_ins_503 : _GEN_502;
  assign _GEN_504 = 9'h1f8 == io_sel ? io_ins_504 : _GEN_503;
  assign _GEN_505 = 9'h1f9 == io_sel ? io_ins_505 : _GEN_504;
  assign io_out = _GEN_0;
  assign _GEN_0 = _GEN_505;
endmodule
module RegFile(
  input         clock,
  input         reset,
  input  [31:0] io_raddr,
  input         io_wen,
  input  [31:0] io_waddr,
  input  [63:0] io_wdata,
  output [63:0] io_rdata,
  input         io_reset,
  output [63:0] io_argIns_0,
  output [63:0] io_argIns_1,
  output [63:0] io_argIns_2,
  output [63:0] io_argIns_3,
  output [63:0] io_argIns_4,
  input         io_argOuts_0_valid,
  input  [63:0] io_argOuts_0_bits,
  input         io_argOuts_1_valid,
  input  [63:0] io_argOuts_1_bits,
  input  [63:0] io_argOuts_2_bits,
  input  [63:0] io_argOuts_3_bits,
  input  [63:0] io_argOuts_4_bits,
  input  [63:0] io_argOuts_5_bits,
  input  [63:0] io_argOuts_6_bits,
  input  [63:0] io_argOuts_7_bits,
  input  [63:0] io_argOuts_8_bits,
  input  [63:0] io_argOuts_9_bits,
  input  [63:0] io_argOuts_10_bits,
  input  [63:0] io_argOuts_11_bits,
  input  [63:0] io_argOuts_12_bits,
  input  [63:0] io_argOuts_13_bits,
  input  [63:0] io_argOuts_14_bits,
  input  [63:0] io_argOuts_15_bits,
  input  [63:0] io_argOuts_16_bits,
  input  [63:0] io_argOuts_17_bits,
  input  [63:0] io_argOuts_18_bits,
  input  [63:0] io_argOuts_19_bits,
  input  [63:0] io_argOuts_20_bits,
  input  [63:0] io_argOuts_21_bits,
  input  [63:0] io_argOuts_22_bits,
  input  [63:0] io_argOuts_23_bits,
  input  [63:0] io_argOuts_24_bits,
  input  [63:0] io_argOuts_25_bits,
  input  [63:0] io_argOuts_26_bits,
  input  [63:0] io_argOuts_27_bits,
  input  [63:0] io_argOuts_28_bits,
  input  [63:0] io_argOuts_29_bits,
  input  [63:0] io_argOuts_30_bits,
  input  [63:0] io_argOuts_31_bits,
  input  [63:0] io_argOuts_32_bits,
  input  [63:0] io_argOuts_33_bits,
  input  [63:0] io_argOuts_34_bits,
  input  [63:0] io_argOuts_35_bits,
  input  [63:0] io_argOuts_36_bits,
  input  [63:0] io_argOuts_37_bits,
  input  [63:0] io_argOuts_38_bits,
  input  [63:0] io_argOuts_39_bits,
  input  [63:0] io_argOuts_40_bits,
  input  [63:0] io_argOuts_41_bits,
  input  [63:0] io_argOuts_42_bits,
  input  [63:0] io_argOuts_43_bits,
  input  [63:0] io_argOuts_44_bits,
  input  [63:0] io_argOuts_45_bits,
  input  [63:0] io_argOuts_46_bits,
  input  [63:0] io_argOuts_47_bits,
  input  [63:0] io_argOuts_48_bits,
  input  [63:0] io_argOuts_49_bits,
  input  [63:0] io_argOuts_50_bits,
  input  [63:0] io_argOuts_51_bits,
  input  [63:0] io_argOuts_52_bits,
  input  [63:0] io_argOuts_53_bits,
  input  [63:0] io_argOuts_54_bits,
  input  [63:0] io_argOuts_55_bits,
  input  [63:0] io_argOuts_56_bits,
  input  [63:0] io_argOuts_57_bits,
  input  [63:0] io_argOuts_58_bits,
  input  [63:0] io_argOuts_59_bits,
  input  [63:0] io_argOuts_60_bits,
  input  [63:0] io_argOuts_61_bits,
  input  [63:0] io_argOuts_62_bits,
  input  [63:0] io_argOuts_63_bits,
  input  [63:0] io_argOuts_64_bits,
  input  [63:0] io_argOuts_65_bits,
  input  [63:0] io_argOuts_66_bits,
  input  [63:0] io_argOuts_67_bits,
  input  [63:0] io_argOuts_68_bits,
  input  [63:0] io_argOuts_69_bits,
  input  [63:0] io_argOuts_70_bits,
  input  [63:0] io_argOuts_71_bits,
  input  [63:0] io_argOuts_72_bits,
  input  [63:0] io_argOuts_73_bits,
  input  [63:0] io_argOuts_74_bits,
  input  [63:0] io_argOuts_75_bits,
  input  [63:0] io_argOuts_76_bits,
  input  [63:0] io_argOuts_77_bits,
  input  [63:0] io_argOuts_78_bits,
  input  [63:0] io_argOuts_79_bits,
  input  [63:0] io_argOuts_80_bits,
  input  [63:0] io_argOuts_81_bits,
  input  [63:0] io_argOuts_82_bits,
  input  [63:0] io_argOuts_83_bits,
  input  [63:0] io_argOuts_84_bits,
  input  [63:0] io_argOuts_85_bits,
  input  [63:0] io_argOuts_86_bits,
  input  [63:0] io_argOuts_87_bits,
  input  [63:0] io_argOuts_88_bits,
  input  [63:0] io_argOuts_89_bits,
  input  [63:0] io_argOuts_90_bits,
  input  [63:0] io_argOuts_91_bits,
  input  [63:0] io_argOuts_92_bits,
  input  [63:0] io_argOuts_93_bits,
  input  [63:0] io_argOuts_94_bits,
  input  [63:0] io_argOuts_95_bits,
  input  [63:0] io_argOuts_96_bits,
  input  [63:0] io_argOuts_97_bits,
  input  [63:0] io_argOuts_98_bits,
  input  [63:0] io_argOuts_99_bits,
  input  [63:0] io_argOuts_100_bits,
  input  [63:0] io_argOuts_101_bits,
  input  [63:0] io_argOuts_102_bits,
  input  [63:0] io_argOuts_103_bits,
  input  [63:0] io_argOuts_104_bits,
  input  [63:0] io_argOuts_105_bits,
  input  [63:0] io_argOuts_106_bits,
  input  [63:0] io_argOuts_107_bits,
  input  [63:0] io_argOuts_108_bits,
  input  [63:0] io_argOuts_109_bits
);
  wire  regs_0_clock;
  wire  regs_0_reset;
  wire [63:0] regs_0_io_in;
  wire [63:0] regs_0_io_init;
  wire  regs_0_io_reset;
  wire [63:0] regs_0_io_out;
  wire  regs_0_io_enable;
  wire  _T_1544;
  wire  _T_1545;
  wire  regs_1_clock;
  wire  regs_1_reset;
  wire [63:0] regs_1_io_in;
  wire [63:0] regs_1_io_init;
  wire  regs_1_io_reset;
  wire [63:0] regs_1_io_out;
  wire  regs_1_io_enable;
  wire  _T_1550;
  wire  _T_1551;
  wire  _T_1555;
  wire [63:0] _T_1559;
  wire  regs_2_clock;
  wire  regs_2_reset;
  wire [63:0] regs_2_io_in;
  wire [63:0] regs_2_io_init;
  wire  regs_2_io_reset;
  wire [63:0] regs_2_io_out;
  wire  regs_2_io_enable;
  wire  _T_1564;
  wire  _T_1565;
  wire  regs_3_clock;
  wire  regs_3_reset;
  wire [63:0] regs_3_io_in;
  wire [63:0] regs_3_io_init;
  wire  regs_3_io_reset;
  wire [63:0] regs_3_io_out;
  wire  regs_3_io_enable;
  wire  _T_1570;
  wire  _T_1571;
  wire  regs_4_clock;
  wire  regs_4_reset;
  wire [63:0] regs_4_io_in;
  wire [63:0] regs_4_io_init;
  wire  regs_4_io_reset;
  wire [63:0] regs_4_io_out;
  wire  regs_4_io_enable;
  wire  _T_1576;
  wire  _T_1577;
  wire  regs_5_clock;
  wire  regs_5_reset;
  wire [63:0] regs_5_io_in;
  wire [63:0] regs_5_io_init;
  wire  regs_5_io_reset;
  wire [63:0] regs_5_io_out;
  wire  regs_5_io_enable;
  wire  _T_1582;
  wire  _T_1583;
  wire  _T_1584;
  wire [63:0] _T_1585;
  wire  regs_6_clock;
  wire  regs_6_reset;
  wire [63:0] regs_6_io_in;
  wire [63:0] regs_6_io_init;
  wire  regs_6_io_reset;
  wire [63:0] regs_6_io_out;
  wire  regs_6_io_enable;
  wire  regs_7_clock;
  wire  regs_7_reset;
  wire [63:0] regs_7_io_in;
  wire [63:0] regs_7_io_init;
  wire  regs_7_io_reset;
  wire [63:0] regs_7_io_out;
  wire  regs_7_io_enable;
  wire  regs_8_clock;
  wire  regs_8_reset;
  wire [63:0] regs_8_io_in;
  wire [63:0] regs_8_io_init;
  wire  regs_8_io_reset;
  wire [63:0] regs_8_io_out;
  wire  regs_8_io_enable;
  wire  regs_9_clock;
  wire  regs_9_reset;
  wire [63:0] regs_9_io_in;
  wire [63:0] regs_9_io_init;
  wire  regs_9_io_reset;
  wire [63:0] regs_9_io_out;
  wire  regs_9_io_enable;
  wire  regs_10_clock;
  wire  regs_10_reset;
  wire [63:0] regs_10_io_in;
  wire [63:0] regs_10_io_init;
  wire  regs_10_io_reset;
  wire [63:0] regs_10_io_out;
  wire  regs_10_io_enable;
  wire  regs_11_clock;
  wire  regs_11_reset;
  wire [63:0] regs_11_io_in;
  wire [63:0] regs_11_io_init;
  wire  regs_11_io_reset;
  wire [63:0] regs_11_io_out;
  wire  regs_11_io_enable;
  wire  regs_12_clock;
  wire  regs_12_reset;
  wire [63:0] regs_12_io_in;
  wire [63:0] regs_12_io_init;
  wire  regs_12_io_reset;
  wire [63:0] regs_12_io_out;
  wire  regs_12_io_enable;
  wire  regs_13_clock;
  wire  regs_13_reset;
  wire [63:0] regs_13_io_in;
  wire [63:0] regs_13_io_init;
  wire  regs_13_io_reset;
  wire [63:0] regs_13_io_out;
  wire  regs_13_io_enable;
  wire  regs_14_clock;
  wire  regs_14_reset;
  wire [63:0] regs_14_io_in;
  wire [63:0] regs_14_io_init;
  wire  regs_14_io_reset;
  wire [63:0] regs_14_io_out;
  wire  regs_14_io_enable;
  wire  regs_15_clock;
  wire  regs_15_reset;
  wire [63:0] regs_15_io_in;
  wire [63:0] regs_15_io_init;
  wire  regs_15_io_reset;
  wire [63:0] regs_15_io_out;
  wire  regs_15_io_enable;
  wire  regs_16_clock;
  wire  regs_16_reset;
  wire [63:0] regs_16_io_in;
  wire [63:0] regs_16_io_init;
  wire  regs_16_io_reset;
  wire [63:0] regs_16_io_out;
  wire  regs_16_io_enable;
  wire  regs_17_clock;
  wire  regs_17_reset;
  wire [63:0] regs_17_io_in;
  wire [63:0] regs_17_io_init;
  wire  regs_17_io_reset;
  wire [63:0] regs_17_io_out;
  wire  regs_17_io_enable;
  wire  regs_18_clock;
  wire  regs_18_reset;
  wire [63:0] regs_18_io_in;
  wire [63:0] regs_18_io_init;
  wire  regs_18_io_reset;
  wire [63:0] regs_18_io_out;
  wire  regs_18_io_enable;
  wire  regs_19_clock;
  wire  regs_19_reset;
  wire [63:0] regs_19_io_in;
  wire [63:0] regs_19_io_init;
  wire  regs_19_io_reset;
  wire [63:0] regs_19_io_out;
  wire  regs_19_io_enable;
  wire  regs_20_clock;
  wire  regs_20_reset;
  wire [63:0] regs_20_io_in;
  wire [63:0] regs_20_io_init;
  wire  regs_20_io_reset;
  wire [63:0] regs_20_io_out;
  wire  regs_20_io_enable;
  wire  regs_21_clock;
  wire  regs_21_reset;
  wire [63:0] regs_21_io_in;
  wire [63:0] regs_21_io_init;
  wire  regs_21_io_reset;
  wire [63:0] regs_21_io_out;
  wire  regs_21_io_enable;
  wire  regs_22_clock;
  wire  regs_22_reset;
  wire [63:0] regs_22_io_in;
  wire [63:0] regs_22_io_init;
  wire  regs_22_io_reset;
  wire [63:0] regs_22_io_out;
  wire  regs_22_io_enable;
  wire  regs_23_clock;
  wire  regs_23_reset;
  wire [63:0] regs_23_io_in;
  wire [63:0] regs_23_io_init;
  wire  regs_23_io_reset;
  wire [63:0] regs_23_io_out;
  wire  regs_23_io_enable;
  wire  regs_24_clock;
  wire  regs_24_reset;
  wire [63:0] regs_24_io_in;
  wire [63:0] regs_24_io_init;
  wire  regs_24_io_reset;
  wire [63:0] regs_24_io_out;
  wire  regs_24_io_enable;
  wire  regs_25_clock;
  wire  regs_25_reset;
  wire [63:0] regs_25_io_in;
  wire [63:0] regs_25_io_init;
  wire  regs_25_io_reset;
  wire [63:0] regs_25_io_out;
  wire  regs_25_io_enable;
  wire  regs_26_clock;
  wire  regs_26_reset;
  wire [63:0] regs_26_io_in;
  wire [63:0] regs_26_io_init;
  wire  regs_26_io_reset;
  wire [63:0] regs_26_io_out;
  wire  regs_26_io_enable;
  wire  regs_27_clock;
  wire  regs_27_reset;
  wire [63:0] regs_27_io_in;
  wire [63:0] regs_27_io_init;
  wire  regs_27_io_reset;
  wire [63:0] regs_27_io_out;
  wire  regs_27_io_enable;
  wire  regs_28_clock;
  wire  regs_28_reset;
  wire [63:0] regs_28_io_in;
  wire [63:0] regs_28_io_init;
  wire  regs_28_io_reset;
  wire [63:0] regs_28_io_out;
  wire  regs_28_io_enable;
  wire  regs_29_clock;
  wire  regs_29_reset;
  wire [63:0] regs_29_io_in;
  wire [63:0] regs_29_io_init;
  wire  regs_29_io_reset;
  wire [63:0] regs_29_io_out;
  wire  regs_29_io_enable;
  wire  regs_30_clock;
  wire  regs_30_reset;
  wire [63:0] regs_30_io_in;
  wire [63:0] regs_30_io_init;
  wire  regs_30_io_reset;
  wire [63:0] regs_30_io_out;
  wire  regs_30_io_enable;
  wire  regs_31_clock;
  wire  regs_31_reset;
  wire [63:0] regs_31_io_in;
  wire [63:0] regs_31_io_init;
  wire  regs_31_io_reset;
  wire [63:0] regs_31_io_out;
  wire  regs_31_io_enable;
  wire  regs_32_clock;
  wire  regs_32_reset;
  wire [63:0] regs_32_io_in;
  wire [63:0] regs_32_io_init;
  wire  regs_32_io_reset;
  wire [63:0] regs_32_io_out;
  wire  regs_32_io_enable;
  wire  regs_33_clock;
  wire  regs_33_reset;
  wire [63:0] regs_33_io_in;
  wire [63:0] regs_33_io_init;
  wire  regs_33_io_reset;
  wire [63:0] regs_33_io_out;
  wire  regs_33_io_enable;
  wire  regs_34_clock;
  wire  regs_34_reset;
  wire [63:0] regs_34_io_in;
  wire [63:0] regs_34_io_init;
  wire  regs_34_io_reset;
  wire [63:0] regs_34_io_out;
  wire  regs_34_io_enable;
  wire  regs_35_clock;
  wire  regs_35_reset;
  wire [63:0] regs_35_io_in;
  wire [63:0] regs_35_io_init;
  wire  regs_35_io_reset;
  wire [63:0] regs_35_io_out;
  wire  regs_35_io_enable;
  wire  regs_36_clock;
  wire  regs_36_reset;
  wire [63:0] regs_36_io_in;
  wire [63:0] regs_36_io_init;
  wire  regs_36_io_reset;
  wire [63:0] regs_36_io_out;
  wire  regs_36_io_enable;
  wire  regs_37_clock;
  wire  regs_37_reset;
  wire [63:0] regs_37_io_in;
  wire [63:0] regs_37_io_init;
  wire  regs_37_io_reset;
  wire [63:0] regs_37_io_out;
  wire  regs_37_io_enable;
  wire  regs_38_clock;
  wire  regs_38_reset;
  wire [63:0] regs_38_io_in;
  wire [63:0] regs_38_io_init;
  wire  regs_38_io_reset;
  wire [63:0] regs_38_io_out;
  wire  regs_38_io_enable;
  wire  regs_39_clock;
  wire  regs_39_reset;
  wire [63:0] regs_39_io_in;
  wire [63:0] regs_39_io_init;
  wire  regs_39_io_reset;
  wire [63:0] regs_39_io_out;
  wire  regs_39_io_enable;
  wire  regs_40_clock;
  wire  regs_40_reset;
  wire [63:0] regs_40_io_in;
  wire [63:0] regs_40_io_init;
  wire  regs_40_io_reset;
  wire [63:0] regs_40_io_out;
  wire  regs_40_io_enable;
  wire  regs_41_clock;
  wire  regs_41_reset;
  wire [63:0] regs_41_io_in;
  wire [63:0] regs_41_io_init;
  wire  regs_41_io_reset;
  wire [63:0] regs_41_io_out;
  wire  regs_41_io_enable;
  wire  regs_42_clock;
  wire  regs_42_reset;
  wire [63:0] regs_42_io_in;
  wire [63:0] regs_42_io_init;
  wire  regs_42_io_reset;
  wire [63:0] regs_42_io_out;
  wire  regs_42_io_enable;
  wire  regs_43_clock;
  wire  regs_43_reset;
  wire [63:0] regs_43_io_in;
  wire [63:0] regs_43_io_init;
  wire  regs_43_io_reset;
  wire [63:0] regs_43_io_out;
  wire  regs_43_io_enable;
  wire  regs_44_clock;
  wire  regs_44_reset;
  wire [63:0] regs_44_io_in;
  wire [63:0] regs_44_io_init;
  wire  regs_44_io_reset;
  wire [63:0] regs_44_io_out;
  wire  regs_44_io_enable;
  wire  regs_45_clock;
  wire  regs_45_reset;
  wire [63:0] regs_45_io_in;
  wire [63:0] regs_45_io_init;
  wire  regs_45_io_reset;
  wire [63:0] regs_45_io_out;
  wire  regs_45_io_enable;
  wire  regs_46_clock;
  wire  regs_46_reset;
  wire [63:0] regs_46_io_in;
  wire [63:0] regs_46_io_init;
  wire  regs_46_io_reset;
  wire [63:0] regs_46_io_out;
  wire  regs_46_io_enable;
  wire  regs_47_clock;
  wire  regs_47_reset;
  wire [63:0] regs_47_io_in;
  wire [63:0] regs_47_io_init;
  wire  regs_47_io_reset;
  wire [63:0] regs_47_io_out;
  wire  regs_47_io_enable;
  wire  regs_48_clock;
  wire  regs_48_reset;
  wire [63:0] regs_48_io_in;
  wire [63:0] regs_48_io_init;
  wire  regs_48_io_reset;
  wire [63:0] regs_48_io_out;
  wire  regs_48_io_enable;
  wire  regs_49_clock;
  wire  regs_49_reset;
  wire [63:0] regs_49_io_in;
  wire [63:0] regs_49_io_init;
  wire  regs_49_io_reset;
  wire [63:0] regs_49_io_out;
  wire  regs_49_io_enable;
  wire  regs_50_clock;
  wire  regs_50_reset;
  wire [63:0] regs_50_io_in;
  wire [63:0] regs_50_io_init;
  wire  regs_50_io_reset;
  wire [63:0] regs_50_io_out;
  wire  regs_50_io_enable;
  wire  regs_51_clock;
  wire  regs_51_reset;
  wire [63:0] regs_51_io_in;
  wire [63:0] regs_51_io_init;
  wire  regs_51_io_reset;
  wire [63:0] regs_51_io_out;
  wire  regs_51_io_enable;
  wire  regs_52_clock;
  wire  regs_52_reset;
  wire [63:0] regs_52_io_in;
  wire [63:0] regs_52_io_init;
  wire  regs_52_io_reset;
  wire [63:0] regs_52_io_out;
  wire  regs_52_io_enable;
  wire  regs_53_clock;
  wire  regs_53_reset;
  wire [63:0] regs_53_io_in;
  wire [63:0] regs_53_io_init;
  wire  regs_53_io_reset;
  wire [63:0] regs_53_io_out;
  wire  regs_53_io_enable;
  wire  regs_54_clock;
  wire  regs_54_reset;
  wire [63:0] regs_54_io_in;
  wire [63:0] regs_54_io_init;
  wire  regs_54_io_reset;
  wire [63:0] regs_54_io_out;
  wire  regs_54_io_enable;
  wire  regs_55_clock;
  wire  regs_55_reset;
  wire [63:0] regs_55_io_in;
  wire [63:0] regs_55_io_init;
  wire  regs_55_io_reset;
  wire [63:0] regs_55_io_out;
  wire  regs_55_io_enable;
  wire  regs_56_clock;
  wire  regs_56_reset;
  wire [63:0] regs_56_io_in;
  wire [63:0] regs_56_io_init;
  wire  regs_56_io_reset;
  wire [63:0] regs_56_io_out;
  wire  regs_56_io_enable;
  wire  regs_57_clock;
  wire  regs_57_reset;
  wire [63:0] regs_57_io_in;
  wire [63:0] regs_57_io_init;
  wire  regs_57_io_reset;
  wire [63:0] regs_57_io_out;
  wire  regs_57_io_enable;
  wire  regs_58_clock;
  wire  regs_58_reset;
  wire [63:0] regs_58_io_in;
  wire [63:0] regs_58_io_init;
  wire  regs_58_io_reset;
  wire [63:0] regs_58_io_out;
  wire  regs_58_io_enable;
  wire  regs_59_clock;
  wire  regs_59_reset;
  wire [63:0] regs_59_io_in;
  wire [63:0] regs_59_io_init;
  wire  regs_59_io_reset;
  wire [63:0] regs_59_io_out;
  wire  regs_59_io_enable;
  wire  regs_60_clock;
  wire  regs_60_reset;
  wire [63:0] regs_60_io_in;
  wire [63:0] regs_60_io_init;
  wire  regs_60_io_reset;
  wire [63:0] regs_60_io_out;
  wire  regs_60_io_enable;
  wire  regs_61_clock;
  wire  regs_61_reset;
  wire [63:0] regs_61_io_in;
  wire [63:0] regs_61_io_init;
  wire  regs_61_io_reset;
  wire [63:0] regs_61_io_out;
  wire  regs_61_io_enable;
  wire  regs_62_clock;
  wire  regs_62_reset;
  wire [63:0] regs_62_io_in;
  wire [63:0] regs_62_io_init;
  wire  regs_62_io_reset;
  wire [63:0] regs_62_io_out;
  wire  regs_62_io_enable;
  wire  regs_63_clock;
  wire  regs_63_reset;
  wire [63:0] regs_63_io_in;
  wire [63:0] regs_63_io_init;
  wire  regs_63_io_reset;
  wire [63:0] regs_63_io_out;
  wire  regs_63_io_enable;
  wire  regs_64_clock;
  wire  regs_64_reset;
  wire [63:0] regs_64_io_in;
  wire [63:0] regs_64_io_init;
  wire  regs_64_io_reset;
  wire [63:0] regs_64_io_out;
  wire  regs_64_io_enable;
  wire  regs_65_clock;
  wire  regs_65_reset;
  wire [63:0] regs_65_io_in;
  wire [63:0] regs_65_io_init;
  wire  regs_65_io_reset;
  wire [63:0] regs_65_io_out;
  wire  regs_65_io_enable;
  wire  regs_66_clock;
  wire  regs_66_reset;
  wire [63:0] regs_66_io_in;
  wire [63:0] regs_66_io_init;
  wire  regs_66_io_reset;
  wire [63:0] regs_66_io_out;
  wire  regs_66_io_enable;
  wire  regs_67_clock;
  wire  regs_67_reset;
  wire [63:0] regs_67_io_in;
  wire [63:0] regs_67_io_init;
  wire  regs_67_io_reset;
  wire [63:0] regs_67_io_out;
  wire  regs_67_io_enable;
  wire  regs_68_clock;
  wire  regs_68_reset;
  wire [63:0] regs_68_io_in;
  wire [63:0] regs_68_io_init;
  wire  regs_68_io_reset;
  wire [63:0] regs_68_io_out;
  wire  regs_68_io_enable;
  wire  regs_69_clock;
  wire  regs_69_reset;
  wire [63:0] regs_69_io_in;
  wire [63:0] regs_69_io_init;
  wire  regs_69_io_reset;
  wire [63:0] regs_69_io_out;
  wire  regs_69_io_enable;
  wire  regs_70_clock;
  wire  regs_70_reset;
  wire [63:0] regs_70_io_in;
  wire [63:0] regs_70_io_init;
  wire  regs_70_io_reset;
  wire [63:0] regs_70_io_out;
  wire  regs_70_io_enable;
  wire  regs_71_clock;
  wire  regs_71_reset;
  wire [63:0] regs_71_io_in;
  wire [63:0] regs_71_io_init;
  wire  regs_71_io_reset;
  wire [63:0] regs_71_io_out;
  wire  regs_71_io_enable;
  wire  regs_72_clock;
  wire  regs_72_reset;
  wire [63:0] regs_72_io_in;
  wire [63:0] regs_72_io_init;
  wire  regs_72_io_reset;
  wire [63:0] regs_72_io_out;
  wire  regs_72_io_enable;
  wire  regs_73_clock;
  wire  regs_73_reset;
  wire [63:0] regs_73_io_in;
  wire [63:0] regs_73_io_init;
  wire  regs_73_io_reset;
  wire [63:0] regs_73_io_out;
  wire  regs_73_io_enable;
  wire  regs_74_clock;
  wire  regs_74_reset;
  wire [63:0] regs_74_io_in;
  wire [63:0] regs_74_io_init;
  wire  regs_74_io_reset;
  wire [63:0] regs_74_io_out;
  wire  regs_74_io_enable;
  wire  regs_75_clock;
  wire  regs_75_reset;
  wire [63:0] regs_75_io_in;
  wire [63:0] regs_75_io_init;
  wire  regs_75_io_reset;
  wire [63:0] regs_75_io_out;
  wire  regs_75_io_enable;
  wire  regs_76_clock;
  wire  regs_76_reset;
  wire [63:0] regs_76_io_in;
  wire [63:0] regs_76_io_init;
  wire  regs_76_io_reset;
  wire [63:0] regs_76_io_out;
  wire  regs_76_io_enable;
  wire  regs_77_clock;
  wire  regs_77_reset;
  wire [63:0] regs_77_io_in;
  wire [63:0] regs_77_io_init;
  wire  regs_77_io_reset;
  wire [63:0] regs_77_io_out;
  wire  regs_77_io_enable;
  wire  regs_78_clock;
  wire  regs_78_reset;
  wire [63:0] regs_78_io_in;
  wire [63:0] regs_78_io_init;
  wire  regs_78_io_reset;
  wire [63:0] regs_78_io_out;
  wire  regs_78_io_enable;
  wire  regs_79_clock;
  wire  regs_79_reset;
  wire [63:0] regs_79_io_in;
  wire [63:0] regs_79_io_init;
  wire  regs_79_io_reset;
  wire [63:0] regs_79_io_out;
  wire  regs_79_io_enable;
  wire  regs_80_clock;
  wire  regs_80_reset;
  wire [63:0] regs_80_io_in;
  wire [63:0] regs_80_io_init;
  wire  regs_80_io_reset;
  wire [63:0] regs_80_io_out;
  wire  regs_80_io_enable;
  wire  regs_81_clock;
  wire  regs_81_reset;
  wire [63:0] regs_81_io_in;
  wire [63:0] regs_81_io_init;
  wire  regs_81_io_reset;
  wire [63:0] regs_81_io_out;
  wire  regs_81_io_enable;
  wire  regs_82_clock;
  wire  regs_82_reset;
  wire [63:0] regs_82_io_in;
  wire [63:0] regs_82_io_init;
  wire  regs_82_io_reset;
  wire [63:0] regs_82_io_out;
  wire  regs_82_io_enable;
  wire  regs_83_clock;
  wire  regs_83_reset;
  wire [63:0] regs_83_io_in;
  wire [63:0] regs_83_io_init;
  wire  regs_83_io_reset;
  wire [63:0] regs_83_io_out;
  wire  regs_83_io_enable;
  wire  regs_84_clock;
  wire  regs_84_reset;
  wire [63:0] regs_84_io_in;
  wire [63:0] regs_84_io_init;
  wire  regs_84_io_reset;
  wire [63:0] regs_84_io_out;
  wire  regs_84_io_enable;
  wire  regs_85_clock;
  wire  regs_85_reset;
  wire [63:0] regs_85_io_in;
  wire [63:0] regs_85_io_init;
  wire  regs_85_io_reset;
  wire [63:0] regs_85_io_out;
  wire  regs_85_io_enable;
  wire  regs_86_clock;
  wire  regs_86_reset;
  wire [63:0] regs_86_io_in;
  wire [63:0] regs_86_io_init;
  wire  regs_86_io_reset;
  wire [63:0] regs_86_io_out;
  wire  regs_86_io_enable;
  wire  regs_87_clock;
  wire  regs_87_reset;
  wire [63:0] regs_87_io_in;
  wire [63:0] regs_87_io_init;
  wire  regs_87_io_reset;
  wire [63:0] regs_87_io_out;
  wire  regs_87_io_enable;
  wire  regs_88_clock;
  wire  regs_88_reset;
  wire [63:0] regs_88_io_in;
  wire [63:0] regs_88_io_init;
  wire  regs_88_io_reset;
  wire [63:0] regs_88_io_out;
  wire  regs_88_io_enable;
  wire  regs_89_clock;
  wire  regs_89_reset;
  wire [63:0] regs_89_io_in;
  wire [63:0] regs_89_io_init;
  wire  regs_89_io_reset;
  wire [63:0] regs_89_io_out;
  wire  regs_89_io_enable;
  wire  regs_90_clock;
  wire  regs_90_reset;
  wire [63:0] regs_90_io_in;
  wire [63:0] regs_90_io_init;
  wire  regs_90_io_reset;
  wire [63:0] regs_90_io_out;
  wire  regs_90_io_enable;
  wire  regs_91_clock;
  wire  regs_91_reset;
  wire [63:0] regs_91_io_in;
  wire [63:0] regs_91_io_init;
  wire  regs_91_io_reset;
  wire [63:0] regs_91_io_out;
  wire  regs_91_io_enable;
  wire  regs_92_clock;
  wire  regs_92_reset;
  wire [63:0] regs_92_io_in;
  wire [63:0] regs_92_io_init;
  wire  regs_92_io_reset;
  wire [63:0] regs_92_io_out;
  wire  regs_92_io_enable;
  wire  regs_93_clock;
  wire  regs_93_reset;
  wire [63:0] regs_93_io_in;
  wire [63:0] regs_93_io_init;
  wire  regs_93_io_reset;
  wire [63:0] regs_93_io_out;
  wire  regs_93_io_enable;
  wire  regs_94_clock;
  wire  regs_94_reset;
  wire [63:0] regs_94_io_in;
  wire [63:0] regs_94_io_init;
  wire  regs_94_io_reset;
  wire [63:0] regs_94_io_out;
  wire  regs_94_io_enable;
  wire  regs_95_clock;
  wire  regs_95_reset;
  wire [63:0] regs_95_io_in;
  wire [63:0] regs_95_io_init;
  wire  regs_95_io_reset;
  wire [63:0] regs_95_io_out;
  wire  regs_95_io_enable;
  wire  regs_96_clock;
  wire  regs_96_reset;
  wire [63:0] regs_96_io_in;
  wire [63:0] regs_96_io_init;
  wire  regs_96_io_reset;
  wire [63:0] regs_96_io_out;
  wire  regs_96_io_enable;
  wire  regs_97_clock;
  wire  regs_97_reset;
  wire [63:0] regs_97_io_in;
  wire [63:0] regs_97_io_init;
  wire  regs_97_io_reset;
  wire [63:0] regs_97_io_out;
  wire  regs_97_io_enable;
  wire  regs_98_clock;
  wire  regs_98_reset;
  wire [63:0] regs_98_io_in;
  wire [63:0] regs_98_io_init;
  wire  regs_98_io_reset;
  wire [63:0] regs_98_io_out;
  wire  regs_98_io_enable;
  wire  regs_99_clock;
  wire  regs_99_reset;
  wire [63:0] regs_99_io_in;
  wire [63:0] regs_99_io_init;
  wire  regs_99_io_reset;
  wire [63:0] regs_99_io_out;
  wire  regs_99_io_enable;
  wire  regs_100_clock;
  wire  regs_100_reset;
  wire [63:0] regs_100_io_in;
  wire [63:0] regs_100_io_init;
  wire  regs_100_io_reset;
  wire [63:0] regs_100_io_out;
  wire  regs_100_io_enable;
  wire  regs_101_clock;
  wire  regs_101_reset;
  wire [63:0] regs_101_io_in;
  wire [63:0] regs_101_io_init;
  wire  regs_101_io_reset;
  wire [63:0] regs_101_io_out;
  wire  regs_101_io_enable;
  wire  regs_102_clock;
  wire  regs_102_reset;
  wire [63:0] regs_102_io_in;
  wire [63:0] regs_102_io_init;
  wire  regs_102_io_reset;
  wire [63:0] regs_102_io_out;
  wire  regs_102_io_enable;
  wire  regs_103_clock;
  wire  regs_103_reset;
  wire [63:0] regs_103_io_in;
  wire [63:0] regs_103_io_init;
  wire  regs_103_io_reset;
  wire [63:0] regs_103_io_out;
  wire  regs_103_io_enable;
  wire  regs_104_clock;
  wire  regs_104_reset;
  wire [63:0] regs_104_io_in;
  wire [63:0] regs_104_io_init;
  wire  regs_104_io_reset;
  wire [63:0] regs_104_io_out;
  wire  regs_104_io_enable;
  wire  regs_105_clock;
  wire  regs_105_reset;
  wire [63:0] regs_105_io_in;
  wire [63:0] regs_105_io_init;
  wire  regs_105_io_reset;
  wire [63:0] regs_105_io_out;
  wire  regs_105_io_enable;
  wire  regs_106_clock;
  wire  regs_106_reset;
  wire [63:0] regs_106_io_in;
  wire [63:0] regs_106_io_init;
  wire  regs_106_io_reset;
  wire [63:0] regs_106_io_out;
  wire  regs_106_io_enable;
  wire  regs_107_clock;
  wire  regs_107_reset;
  wire [63:0] regs_107_io_in;
  wire [63:0] regs_107_io_init;
  wire  regs_107_io_reset;
  wire [63:0] regs_107_io_out;
  wire  regs_107_io_enable;
  wire  regs_108_clock;
  wire  regs_108_reset;
  wire [63:0] regs_108_io_in;
  wire [63:0] regs_108_io_init;
  wire  regs_108_io_reset;
  wire [63:0] regs_108_io_out;
  wire  regs_108_io_enable;
  wire  regs_109_clock;
  wire  regs_109_reset;
  wire [63:0] regs_109_io_in;
  wire [63:0] regs_109_io_init;
  wire  regs_109_io_reset;
  wire [63:0] regs_109_io_out;
  wire  regs_109_io_enable;
  wire  regs_110_clock;
  wire  regs_110_reset;
  wire [63:0] regs_110_io_in;
  wire [63:0] regs_110_io_init;
  wire  regs_110_io_reset;
  wire [63:0] regs_110_io_out;
  wire  regs_110_io_enable;
  wire  regs_111_clock;
  wire  regs_111_reset;
  wire [63:0] regs_111_io_in;
  wire [63:0] regs_111_io_init;
  wire  regs_111_io_reset;
  wire [63:0] regs_111_io_out;
  wire  regs_111_io_enable;
  wire  regs_112_clock;
  wire  regs_112_reset;
  wire [63:0] regs_112_io_in;
  wire [63:0] regs_112_io_init;
  wire  regs_112_io_reset;
  wire [63:0] regs_112_io_out;
  wire  regs_112_io_enable;
  wire  regs_113_clock;
  wire  regs_113_reset;
  wire [63:0] regs_113_io_in;
  wire [63:0] regs_113_io_init;
  wire  regs_113_io_reset;
  wire [63:0] regs_113_io_out;
  wire  regs_113_io_enable;
  wire  regs_114_clock;
  wire  regs_114_reset;
  wire [63:0] regs_114_io_in;
  wire [63:0] regs_114_io_init;
  wire  regs_114_io_reset;
  wire [63:0] regs_114_io_out;
  wire  regs_114_io_enable;
  wire  regs_115_clock;
  wire  regs_115_reset;
  wire [63:0] regs_115_io_in;
  wire [63:0] regs_115_io_init;
  wire  regs_115_io_reset;
  wire [63:0] regs_115_io_out;
  wire  regs_115_io_enable;
  wire  regs_116_clock;
  wire  regs_116_reset;
  wire [63:0] regs_116_io_in;
  wire [63:0] regs_116_io_init;
  wire  regs_116_io_reset;
  wire [63:0] regs_116_io_out;
  wire  regs_116_io_enable;
  wire  regs_117_clock;
  wire  regs_117_reset;
  wire [63:0] regs_117_io_in;
  wire [63:0] regs_117_io_init;
  wire  regs_117_io_reset;
  wire [63:0] regs_117_io_out;
  wire  regs_117_io_enable;
  wire  regs_118_clock;
  wire  regs_118_reset;
  wire [63:0] regs_118_io_in;
  wire [63:0] regs_118_io_init;
  wire  regs_118_io_reset;
  wire [63:0] regs_118_io_out;
  wire  regs_118_io_enable;
  wire  regs_119_clock;
  wire  regs_119_reset;
  wire [63:0] regs_119_io_in;
  wire [63:0] regs_119_io_init;
  wire  regs_119_io_reset;
  wire [63:0] regs_119_io_out;
  wire  regs_119_io_enable;
  wire  regs_120_clock;
  wire  regs_120_reset;
  wire [63:0] regs_120_io_in;
  wire [63:0] regs_120_io_init;
  wire  regs_120_io_reset;
  wire [63:0] regs_120_io_out;
  wire  regs_120_io_enable;
  wire  regs_121_clock;
  wire  regs_121_reset;
  wire [63:0] regs_121_io_in;
  wire [63:0] regs_121_io_init;
  wire  regs_121_io_reset;
  wire [63:0] regs_121_io_out;
  wire  regs_121_io_enable;
  wire  regs_122_clock;
  wire  regs_122_reset;
  wire [63:0] regs_122_io_in;
  wire [63:0] regs_122_io_init;
  wire  regs_122_io_reset;
  wire [63:0] regs_122_io_out;
  wire  regs_122_io_enable;
  wire  regs_123_clock;
  wire  regs_123_reset;
  wire [63:0] regs_123_io_in;
  wire [63:0] regs_123_io_init;
  wire  regs_123_io_reset;
  wire [63:0] regs_123_io_out;
  wire  regs_123_io_enable;
  wire  regs_124_clock;
  wire  regs_124_reset;
  wire [63:0] regs_124_io_in;
  wire [63:0] regs_124_io_init;
  wire  regs_124_io_reset;
  wire [63:0] regs_124_io_out;
  wire  regs_124_io_enable;
  wire  regs_125_clock;
  wire  regs_125_reset;
  wire [63:0] regs_125_io_in;
  wire [63:0] regs_125_io_init;
  wire  regs_125_io_reset;
  wire [63:0] regs_125_io_out;
  wire  regs_125_io_enable;
  wire  regs_126_clock;
  wire  regs_126_reset;
  wire [63:0] regs_126_io_in;
  wire [63:0] regs_126_io_init;
  wire  regs_126_io_reset;
  wire [63:0] regs_126_io_out;
  wire  regs_126_io_enable;
  wire  regs_127_clock;
  wire  regs_127_reset;
  wire [63:0] regs_127_io_in;
  wire [63:0] regs_127_io_init;
  wire  regs_127_io_reset;
  wire [63:0] regs_127_io_out;
  wire  regs_127_io_enable;
  wire  regs_128_clock;
  wire  regs_128_reset;
  wire [63:0] regs_128_io_in;
  wire [63:0] regs_128_io_init;
  wire  regs_128_io_reset;
  wire [63:0] regs_128_io_out;
  wire  regs_128_io_enable;
  wire  regs_129_clock;
  wire  regs_129_reset;
  wire [63:0] regs_129_io_in;
  wire [63:0] regs_129_io_init;
  wire  regs_129_io_reset;
  wire [63:0] regs_129_io_out;
  wire  regs_129_io_enable;
  wire  regs_130_clock;
  wire  regs_130_reset;
  wire [63:0] regs_130_io_in;
  wire [63:0] regs_130_io_init;
  wire  regs_130_io_reset;
  wire [63:0] regs_130_io_out;
  wire  regs_130_io_enable;
  wire  regs_131_clock;
  wire  regs_131_reset;
  wire [63:0] regs_131_io_in;
  wire [63:0] regs_131_io_init;
  wire  regs_131_io_reset;
  wire [63:0] regs_131_io_out;
  wire  regs_131_io_enable;
  wire  regs_132_clock;
  wire  regs_132_reset;
  wire [63:0] regs_132_io_in;
  wire [63:0] regs_132_io_init;
  wire  regs_132_io_reset;
  wire [63:0] regs_132_io_out;
  wire  regs_132_io_enable;
  wire  regs_133_clock;
  wire  regs_133_reset;
  wire [63:0] regs_133_io_in;
  wire [63:0] regs_133_io_init;
  wire  regs_133_io_reset;
  wire [63:0] regs_133_io_out;
  wire  regs_133_io_enable;
  wire  regs_134_clock;
  wire  regs_134_reset;
  wire [63:0] regs_134_io_in;
  wire [63:0] regs_134_io_init;
  wire  regs_134_io_reset;
  wire [63:0] regs_134_io_out;
  wire  regs_134_io_enable;
  wire  regs_135_clock;
  wire  regs_135_reset;
  wire [63:0] regs_135_io_in;
  wire [63:0] regs_135_io_init;
  wire  regs_135_io_reset;
  wire [63:0] regs_135_io_out;
  wire  regs_135_io_enable;
  wire  regs_136_clock;
  wire  regs_136_reset;
  wire [63:0] regs_136_io_in;
  wire [63:0] regs_136_io_init;
  wire  regs_136_io_reset;
  wire [63:0] regs_136_io_out;
  wire  regs_136_io_enable;
  wire  regs_137_clock;
  wire  regs_137_reset;
  wire [63:0] regs_137_io_in;
  wire [63:0] regs_137_io_init;
  wire  regs_137_io_reset;
  wire [63:0] regs_137_io_out;
  wire  regs_137_io_enable;
  wire  regs_138_clock;
  wire  regs_138_reset;
  wire [63:0] regs_138_io_in;
  wire [63:0] regs_138_io_init;
  wire  regs_138_io_reset;
  wire [63:0] regs_138_io_out;
  wire  regs_138_io_enable;
  wire  regs_139_clock;
  wire  regs_139_reset;
  wire [63:0] regs_139_io_in;
  wire [63:0] regs_139_io_init;
  wire  regs_139_io_reset;
  wire [63:0] regs_139_io_out;
  wire  regs_139_io_enable;
  wire  regs_140_clock;
  wire  regs_140_reset;
  wire [63:0] regs_140_io_in;
  wire [63:0] regs_140_io_init;
  wire  regs_140_io_reset;
  wire [63:0] regs_140_io_out;
  wire  regs_140_io_enable;
  wire  regs_141_clock;
  wire  regs_141_reset;
  wire [63:0] regs_141_io_in;
  wire [63:0] regs_141_io_init;
  wire  regs_141_io_reset;
  wire [63:0] regs_141_io_out;
  wire  regs_141_io_enable;
  wire  regs_142_clock;
  wire  regs_142_reset;
  wire [63:0] regs_142_io_in;
  wire [63:0] regs_142_io_init;
  wire  regs_142_io_reset;
  wire [63:0] regs_142_io_out;
  wire  regs_142_io_enable;
  wire  regs_143_clock;
  wire  regs_143_reset;
  wire [63:0] regs_143_io_in;
  wire [63:0] regs_143_io_init;
  wire  regs_143_io_reset;
  wire [63:0] regs_143_io_out;
  wire  regs_143_io_enable;
  wire  regs_144_clock;
  wire  regs_144_reset;
  wire [63:0] regs_144_io_in;
  wire [63:0] regs_144_io_init;
  wire  regs_144_io_reset;
  wire [63:0] regs_144_io_out;
  wire  regs_144_io_enable;
  wire  regs_145_clock;
  wire  regs_145_reset;
  wire [63:0] regs_145_io_in;
  wire [63:0] regs_145_io_init;
  wire  regs_145_io_reset;
  wire [63:0] regs_145_io_out;
  wire  regs_145_io_enable;
  wire  regs_146_clock;
  wire  regs_146_reset;
  wire [63:0] regs_146_io_in;
  wire [63:0] regs_146_io_init;
  wire  regs_146_io_reset;
  wire [63:0] regs_146_io_out;
  wire  regs_146_io_enable;
  wire  regs_147_clock;
  wire  regs_147_reset;
  wire [63:0] regs_147_io_in;
  wire [63:0] regs_147_io_init;
  wire  regs_147_io_reset;
  wire [63:0] regs_147_io_out;
  wire  regs_147_io_enable;
  wire  regs_148_clock;
  wire  regs_148_reset;
  wire [63:0] regs_148_io_in;
  wire [63:0] regs_148_io_init;
  wire  regs_148_io_reset;
  wire [63:0] regs_148_io_out;
  wire  regs_148_io_enable;
  wire  regs_149_clock;
  wire  regs_149_reset;
  wire [63:0] regs_149_io_in;
  wire [63:0] regs_149_io_init;
  wire  regs_149_io_reset;
  wire [63:0] regs_149_io_out;
  wire  regs_149_io_enable;
  wire  regs_150_clock;
  wire  regs_150_reset;
  wire [63:0] regs_150_io_in;
  wire [63:0] regs_150_io_init;
  wire  regs_150_io_reset;
  wire [63:0] regs_150_io_out;
  wire  regs_150_io_enable;
  wire  regs_151_clock;
  wire  regs_151_reset;
  wire [63:0] regs_151_io_in;
  wire [63:0] regs_151_io_init;
  wire  regs_151_io_reset;
  wire [63:0] regs_151_io_out;
  wire  regs_151_io_enable;
  wire  regs_152_clock;
  wire  regs_152_reset;
  wire [63:0] regs_152_io_in;
  wire [63:0] regs_152_io_init;
  wire  regs_152_io_reset;
  wire [63:0] regs_152_io_out;
  wire  regs_152_io_enable;
  wire  regs_153_clock;
  wire  regs_153_reset;
  wire [63:0] regs_153_io_in;
  wire [63:0] regs_153_io_init;
  wire  regs_153_io_reset;
  wire [63:0] regs_153_io_out;
  wire  regs_153_io_enable;
  wire  regs_154_clock;
  wire  regs_154_reset;
  wire [63:0] regs_154_io_in;
  wire [63:0] regs_154_io_init;
  wire  regs_154_io_reset;
  wire [63:0] regs_154_io_out;
  wire  regs_154_io_enable;
  wire  regs_155_clock;
  wire  regs_155_reset;
  wire [63:0] regs_155_io_in;
  wire [63:0] regs_155_io_init;
  wire  regs_155_io_reset;
  wire [63:0] regs_155_io_out;
  wire  regs_155_io_enable;
  wire  regs_156_clock;
  wire  regs_156_reset;
  wire [63:0] regs_156_io_in;
  wire [63:0] regs_156_io_init;
  wire  regs_156_io_reset;
  wire [63:0] regs_156_io_out;
  wire  regs_156_io_enable;
  wire  regs_157_clock;
  wire  regs_157_reset;
  wire [63:0] regs_157_io_in;
  wire [63:0] regs_157_io_init;
  wire  regs_157_io_reset;
  wire [63:0] regs_157_io_out;
  wire  regs_157_io_enable;
  wire  regs_158_clock;
  wire  regs_158_reset;
  wire [63:0] regs_158_io_in;
  wire [63:0] regs_158_io_init;
  wire  regs_158_io_reset;
  wire [63:0] regs_158_io_out;
  wire  regs_158_io_enable;
  wire  regs_159_clock;
  wire  regs_159_reset;
  wire [63:0] regs_159_io_in;
  wire [63:0] regs_159_io_init;
  wire  regs_159_io_reset;
  wire [63:0] regs_159_io_out;
  wire  regs_159_io_enable;
  wire  regs_160_clock;
  wire  regs_160_reset;
  wire [63:0] regs_160_io_in;
  wire [63:0] regs_160_io_init;
  wire  regs_160_io_reset;
  wire [63:0] regs_160_io_out;
  wire  regs_160_io_enable;
  wire  regs_161_clock;
  wire  regs_161_reset;
  wire [63:0] regs_161_io_in;
  wire [63:0] regs_161_io_init;
  wire  regs_161_io_reset;
  wire [63:0] regs_161_io_out;
  wire  regs_161_io_enable;
  wire  regs_162_clock;
  wire  regs_162_reset;
  wire [63:0] regs_162_io_in;
  wire [63:0] regs_162_io_init;
  wire  regs_162_io_reset;
  wire [63:0] regs_162_io_out;
  wire  regs_162_io_enable;
  wire  regs_163_clock;
  wire  regs_163_reset;
  wire [63:0] regs_163_io_in;
  wire [63:0] regs_163_io_init;
  wire  regs_163_io_reset;
  wire [63:0] regs_163_io_out;
  wire  regs_163_io_enable;
  wire  regs_164_clock;
  wire  regs_164_reset;
  wire [63:0] regs_164_io_in;
  wire [63:0] regs_164_io_init;
  wire  regs_164_io_reset;
  wire [63:0] regs_164_io_out;
  wire  regs_164_io_enable;
  wire  regs_165_clock;
  wire  regs_165_reset;
  wire [63:0] regs_165_io_in;
  wire [63:0] regs_165_io_init;
  wire  regs_165_io_reset;
  wire [63:0] regs_165_io_out;
  wire  regs_165_io_enable;
  wire  regs_166_clock;
  wire  regs_166_reset;
  wire [63:0] regs_166_io_in;
  wire [63:0] regs_166_io_init;
  wire  regs_166_io_reset;
  wire [63:0] regs_166_io_out;
  wire  regs_166_io_enable;
  wire  regs_167_clock;
  wire  regs_167_reset;
  wire [63:0] regs_167_io_in;
  wire [63:0] regs_167_io_init;
  wire  regs_167_io_reset;
  wire [63:0] regs_167_io_out;
  wire  regs_167_io_enable;
  wire  regs_168_clock;
  wire  regs_168_reset;
  wire [63:0] regs_168_io_in;
  wire [63:0] regs_168_io_init;
  wire  regs_168_io_reset;
  wire [63:0] regs_168_io_out;
  wire  regs_168_io_enable;
  wire  regs_169_clock;
  wire  regs_169_reset;
  wire [63:0] regs_169_io_in;
  wire [63:0] regs_169_io_init;
  wire  regs_169_io_reset;
  wire [63:0] regs_169_io_out;
  wire  regs_169_io_enable;
  wire  regs_170_clock;
  wire  regs_170_reset;
  wire [63:0] regs_170_io_in;
  wire [63:0] regs_170_io_init;
  wire  regs_170_io_reset;
  wire [63:0] regs_170_io_out;
  wire  regs_170_io_enable;
  wire  regs_171_clock;
  wire  regs_171_reset;
  wire [63:0] regs_171_io_in;
  wire [63:0] regs_171_io_init;
  wire  regs_171_io_reset;
  wire [63:0] regs_171_io_out;
  wire  regs_171_io_enable;
  wire  regs_172_clock;
  wire  regs_172_reset;
  wire [63:0] regs_172_io_in;
  wire [63:0] regs_172_io_init;
  wire  regs_172_io_reset;
  wire [63:0] regs_172_io_out;
  wire  regs_172_io_enable;
  wire  regs_173_clock;
  wire  regs_173_reset;
  wire [63:0] regs_173_io_in;
  wire [63:0] regs_173_io_init;
  wire  regs_173_io_reset;
  wire [63:0] regs_173_io_out;
  wire  regs_173_io_enable;
  wire  regs_174_clock;
  wire  regs_174_reset;
  wire [63:0] regs_174_io_in;
  wire [63:0] regs_174_io_init;
  wire  regs_174_io_reset;
  wire [63:0] regs_174_io_out;
  wire  regs_174_io_enable;
  wire  regs_175_clock;
  wire  regs_175_reset;
  wire [63:0] regs_175_io_in;
  wire [63:0] regs_175_io_init;
  wire  regs_175_io_reset;
  wire [63:0] regs_175_io_out;
  wire  regs_175_io_enable;
  wire  regs_176_clock;
  wire  regs_176_reset;
  wire [63:0] regs_176_io_in;
  wire [63:0] regs_176_io_init;
  wire  regs_176_io_reset;
  wire [63:0] regs_176_io_out;
  wire  regs_176_io_enable;
  wire  regs_177_clock;
  wire  regs_177_reset;
  wire [63:0] regs_177_io_in;
  wire [63:0] regs_177_io_init;
  wire  regs_177_io_reset;
  wire [63:0] regs_177_io_out;
  wire  regs_177_io_enable;
  wire  regs_178_clock;
  wire  regs_178_reset;
  wire [63:0] regs_178_io_in;
  wire [63:0] regs_178_io_init;
  wire  regs_178_io_reset;
  wire [63:0] regs_178_io_out;
  wire  regs_178_io_enable;
  wire  regs_179_clock;
  wire  regs_179_reset;
  wire [63:0] regs_179_io_in;
  wire [63:0] regs_179_io_init;
  wire  regs_179_io_reset;
  wire [63:0] regs_179_io_out;
  wire  regs_179_io_enable;
  wire  regs_180_clock;
  wire  regs_180_reset;
  wire [63:0] regs_180_io_in;
  wire [63:0] regs_180_io_init;
  wire  regs_180_io_reset;
  wire [63:0] regs_180_io_out;
  wire  regs_180_io_enable;
  wire  regs_181_clock;
  wire  regs_181_reset;
  wire [63:0] regs_181_io_in;
  wire [63:0] regs_181_io_init;
  wire  regs_181_io_reset;
  wire [63:0] regs_181_io_out;
  wire  regs_181_io_enable;
  wire  regs_182_clock;
  wire  regs_182_reset;
  wire [63:0] regs_182_io_in;
  wire [63:0] regs_182_io_init;
  wire  regs_182_io_reset;
  wire [63:0] regs_182_io_out;
  wire  regs_182_io_enable;
  wire  regs_183_clock;
  wire  regs_183_reset;
  wire [63:0] regs_183_io_in;
  wire [63:0] regs_183_io_init;
  wire  regs_183_io_reset;
  wire [63:0] regs_183_io_out;
  wire  regs_183_io_enable;
  wire  regs_184_clock;
  wire  regs_184_reset;
  wire [63:0] regs_184_io_in;
  wire [63:0] regs_184_io_init;
  wire  regs_184_io_reset;
  wire [63:0] regs_184_io_out;
  wire  regs_184_io_enable;
  wire  regs_185_clock;
  wire  regs_185_reset;
  wire [63:0] regs_185_io_in;
  wire [63:0] regs_185_io_init;
  wire  regs_185_io_reset;
  wire [63:0] regs_185_io_out;
  wire  regs_185_io_enable;
  wire  regs_186_clock;
  wire  regs_186_reset;
  wire [63:0] regs_186_io_in;
  wire [63:0] regs_186_io_init;
  wire  regs_186_io_reset;
  wire [63:0] regs_186_io_out;
  wire  regs_186_io_enable;
  wire  regs_187_clock;
  wire  regs_187_reset;
  wire [63:0] regs_187_io_in;
  wire [63:0] regs_187_io_init;
  wire  regs_187_io_reset;
  wire [63:0] regs_187_io_out;
  wire  regs_187_io_enable;
  wire  regs_188_clock;
  wire  regs_188_reset;
  wire [63:0] regs_188_io_in;
  wire [63:0] regs_188_io_init;
  wire  regs_188_io_reset;
  wire [63:0] regs_188_io_out;
  wire  regs_188_io_enable;
  wire  regs_189_clock;
  wire  regs_189_reset;
  wire [63:0] regs_189_io_in;
  wire [63:0] regs_189_io_init;
  wire  regs_189_io_reset;
  wire [63:0] regs_189_io_out;
  wire  regs_189_io_enable;
  wire  regs_190_clock;
  wire  regs_190_reset;
  wire [63:0] regs_190_io_in;
  wire [63:0] regs_190_io_init;
  wire  regs_190_io_reset;
  wire [63:0] regs_190_io_out;
  wire  regs_190_io_enable;
  wire  regs_191_clock;
  wire  regs_191_reset;
  wire [63:0] regs_191_io_in;
  wire [63:0] regs_191_io_init;
  wire  regs_191_io_reset;
  wire [63:0] regs_191_io_out;
  wire  regs_191_io_enable;
  wire  regs_192_clock;
  wire  regs_192_reset;
  wire [63:0] regs_192_io_in;
  wire [63:0] regs_192_io_init;
  wire  regs_192_io_reset;
  wire [63:0] regs_192_io_out;
  wire  regs_192_io_enable;
  wire  regs_193_clock;
  wire  regs_193_reset;
  wire [63:0] regs_193_io_in;
  wire [63:0] regs_193_io_init;
  wire  regs_193_io_reset;
  wire [63:0] regs_193_io_out;
  wire  regs_193_io_enable;
  wire  regs_194_clock;
  wire  regs_194_reset;
  wire [63:0] regs_194_io_in;
  wire [63:0] regs_194_io_init;
  wire  regs_194_io_reset;
  wire [63:0] regs_194_io_out;
  wire  regs_194_io_enable;
  wire  regs_195_clock;
  wire  regs_195_reset;
  wire [63:0] regs_195_io_in;
  wire [63:0] regs_195_io_init;
  wire  regs_195_io_reset;
  wire [63:0] regs_195_io_out;
  wire  regs_195_io_enable;
  wire  regs_196_clock;
  wire  regs_196_reset;
  wire [63:0] regs_196_io_in;
  wire [63:0] regs_196_io_init;
  wire  regs_196_io_reset;
  wire [63:0] regs_196_io_out;
  wire  regs_196_io_enable;
  wire  regs_197_clock;
  wire  regs_197_reset;
  wire [63:0] regs_197_io_in;
  wire [63:0] regs_197_io_init;
  wire  regs_197_io_reset;
  wire [63:0] regs_197_io_out;
  wire  regs_197_io_enable;
  wire  regs_198_clock;
  wire  regs_198_reset;
  wire [63:0] regs_198_io_in;
  wire [63:0] regs_198_io_init;
  wire  regs_198_io_reset;
  wire [63:0] regs_198_io_out;
  wire  regs_198_io_enable;
  wire  regs_199_clock;
  wire  regs_199_reset;
  wire [63:0] regs_199_io_in;
  wire [63:0] regs_199_io_init;
  wire  regs_199_io_reset;
  wire [63:0] regs_199_io_out;
  wire  regs_199_io_enable;
  wire  regs_200_clock;
  wire  regs_200_reset;
  wire [63:0] regs_200_io_in;
  wire [63:0] regs_200_io_init;
  wire  regs_200_io_reset;
  wire [63:0] regs_200_io_out;
  wire  regs_200_io_enable;
  wire  regs_201_clock;
  wire  regs_201_reset;
  wire [63:0] regs_201_io_in;
  wire [63:0] regs_201_io_init;
  wire  regs_201_io_reset;
  wire [63:0] regs_201_io_out;
  wire  regs_201_io_enable;
  wire  regs_202_clock;
  wire  regs_202_reset;
  wire [63:0] regs_202_io_in;
  wire [63:0] regs_202_io_init;
  wire  regs_202_io_reset;
  wire [63:0] regs_202_io_out;
  wire  regs_202_io_enable;
  wire  regs_203_clock;
  wire  regs_203_reset;
  wire [63:0] regs_203_io_in;
  wire [63:0] regs_203_io_init;
  wire  regs_203_io_reset;
  wire [63:0] regs_203_io_out;
  wire  regs_203_io_enable;
  wire  regs_204_clock;
  wire  regs_204_reset;
  wire [63:0] regs_204_io_in;
  wire [63:0] regs_204_io_init;
  wire  regs_204_io_reset;
  wire [63:0] regs_204_io_out;
  wire  regs_204_io_enable;
  wire  regs_205_clock;
  wire  regs_205_reset;
  wire [63:0] regs_205_io_in;
  wire [63:0] regs_205_io_init;
  wire  regs_205_io_reset;
  wire [63:0] regs_205_io_out;
  wire  regs_205_io_enable;
  wire  regs_206_clock;
  wire  regs_206_reset;
  wire [63:0] regs_206_io_in;
  wire [63:0] regs_206_io_init;
  wire  regs_206_io_reset;
  wire [63:0] regs_206_io_out;
  wire  regs_206_io_enable;
  wire  regs_207_clock;
  wire  regs_207_reset;
  wire [63:0] regs_207_io_in;
  wire [63:0] regs_207_io_init;
  wire  regs_207_io_reset;
  wire [63:0] regs_207_io_out;
  wire  regs_207_io_enable;
  wire  regs_208_clock;
  wire  regs_208_reset;
  wire [63:0] regs_208_io_in;
  wire [63:0] regs_208_io_init;
  wire  regs_208_io_reset;
  wire [63:0] regs_208_io_out;
  wire  regs_208_io_enable;
  wire  regs_209_clock;
  wire  regs_209_reset;
  wire [63:0] regs_209_io_in;
  wire [63:0] regs_209_io_init;
  wire  regs_209_io_reset;
  wire [63:0] regs_209_io_out;
  wire  regs_209_io_enable;
  wire  regs_210_clock;
  wire  regs_210_reset;
  wire [63:0] regs_210_io_in;
  wire [63:0] regs_210_io_init;
  wire  regs_210_io_reset;
  wire [63:0] regs_210_io_out;
  wire  regs_210_io_enable;
  wire  regs_211_clock;
  wire  regs_211_reset;
  wire [63:0] regs_211_io_in;
  wire [63:0] regs_211_io_init;
  wire  regs_211_io_reset;
  wire [63:0] regs_211_io_out;
  wire  regs_211_io_enable;
  wire  regs_212_clock;
  wire  regs_212_reset;
  wire [63:0] regs_212_io_in;
  wire [63:0] regs_212_io_init;
  wire  regs_212_io_reset;
  wire [63:0] regs_212_io_out;
  wire  regs_212_io_enable;
  wire  regs_213_clock;
  wire  regs_213_reset;
  wire [63:0] regs_213_io_in;
  wire [63:0] regs_213_io_init;
  wire  regs_213_io_reset;
  wire [63:0] regs_213_io_out;
  wire  regs_213_io_enable;
  wire  regs_214_clock;
  wire  regs_214_reset;
  wire [63:0] regs_214_io_in;
  wire [63:0] regs_214_io_init;
  wire  regs_214_io_reset;
  wire [63:0] regs_214_io_out;
  wire  regs_214_io_enable;
  wire  regs_215_clock;
  wire  regs_215_reset;
  wire [63:0] regs_215_io_in;
  wire [63:0] regs_215_io_init;
  wire  regs_215_io_reset;
  wire [63:0] regs_215_io_out;
  wire  regs_215_io_enable;
  wire  regs_216_clock;
  wire  regs_216_reset;
  wire [63:0] regs_216_io_in;
  wire [63:0] regs_216_io_init;
  wire  regs_216_io_reset;
  wire [63:0] regs_216_io_out;
  wire  regs_216_io_enable;
  wire  regs_217_clock;
  wire  regs_217_reset;
  wire [63:0] regs_217_io_in;
  wire [63:0] regs_217_io_init;
  wire  regs_217_io_reset;
  wire [63:0] regs_217_io_out;
  wire  regs_217_io_enable;
  wire  regs_218_clock;
  wire  regs_218_reset;
  wire [63:0] regs_218_io_in;
  wire [63:0] regs_218_io_init;
  wire  regs_218_io_reset;
  wire [63:0] regs_218_io_out;
  wire  regs_218_io_enable;
  wire  regs_219_clock;
  wire  regs_219_reset;
  wire [63:0] regs_219_io_in;
  wire [63:0] regs_219_io_init;
  wire  regs_219_io_reset;
  wire [63:0] regs_219_io_out;
  wire  regs_219_io_enable;
  wire  regs_220_clock;
  wire  regs_220_reset;
  wire [63:0] regs_220_io_in;
  wire [63:0] regs_220_io_init;
  wire  regs_220_io_reset;
  wire [63:0] regs_220_io_out;
  wire  regs_220_io_enable;
  wire  regs_221_clock;
  wire  regs_221_reset;
  wire [63:0] regs_221_io_in;
  wire [63:0] regs_221_io_init;
  wire  regs_221_io_reset;
  wire [63:0] regs_221_io_out;
  wire  regs_221_io_enable;
  wire  regs_222_clock;
  wire  regs_222_reset;
  wire [63:0] regs_222_io_in;
  wire [63:0] regs_222_io_init;
  wire  regs_222_io_reset;
  wire [63:0] regs_222_io_out;
  wire  regs_222_io_enable;
  wire  regs_223_clock;
  wire  regs_223_reset;
  wire [63:0] regs_223_io_in;
  wire [63:0] regs_223_io_init;
  wire  regs_223_io_reset;
  wire [63:0] regs_223_io_out;
  wire  regs_223_io_enable;
  wire  regs_224_clock;
  wire  regs_224_reset;
  wire [63:0] regs_224_io_in;
  wire [63:0] regs_224_io_init;
  wire  regs_224_io_reset;
  wire [63:0] regs_224_io_out;
  wire  regs_224_io_enable;
  wire  regs_225_clock;
  wire  regs_225_reset;
  wire [63:0] regs_225_io_in;
  wire [63:0] regs_225_io_init;
  wire  regs_225_io_reset;
  wire [63:0] regs_225_io_out;
  wire  regs_225_io_enable;
  wire  regs_226_clock;
  wire  regs_226_reset;
  wire [63:0] regs_226_io_in;
  wire [63:0] regs_226_io_init;
  wire  regs_226_io_reset;
  wire [63:0] regs_226_io_out;
  wire  regs_226_io_enable;
  wire  regs_227_clock;
  wire  regs_227_reset;
  wire [63:0] regs_227_io_in;
  wire [63:0] regs_227_io_init;
  wire  regs_227_io_reset;
  wire [63:0] regs_227_io_out;
  wire  regs_227_io_enable;
  wire  regs_228_clock;
  wire  regs_228_reset;
  wire [63:0] regs_228_io_in;
  wire [63:0] regs_228_io_init;
  wire  regs_228_io_reset;
  wire [63:0] regs_228_io_out;
  wire  regs_228_io_enable;
  wire  regs_229_clock;
  wire  regs_229_reset;
  wire [63:0] regs_229_io_in;
  wire [63:0] regs_229_io_init;
  wire  regs_229_io_reset;
  wire [63:0] regs_229_io_out;
  wire  regs_229_io_enable;
  wire  regs_230_clock;
  wire  regs_230_reset;
  wire [63:0] regs_230_io_in;
  wire [63:0] regs_230_io_init;
  wire  regs_230_io_reset;
  wire [63:0] regs_230_io_out;
  wire  regs_230_io_enable;
  wire  regs_231_clock;
  wire  regs_231_reset;
  wire [63:0] regs_231_io_in;
  wire [63:0] regs_231_io_init;
  wire  regs_231_io_reset;
  wire [63:0] regs_231_io_out;
  wire  regs_231_io_enable;
  wire  regs_232_clock;
  wire  regs_232_reset;
  wire [63:0] regs_232_io_in;
  wire [63:0] regs_232_io_init;
  wire  regs_232_io_reset;
  wire [63:0] regs_232_io_out;
  wire  regs_232_io_enable;
  wire  regs_233_clock;
  wire  regs_233_reset;
  wire [63:0] regs_233_io_in;
  wire [63:0] regs_233_io_init;
  wire  regs_233_io_reset;
  wire [63:0] regs_233_io_out;
  wire  regs_233_io_enable;
  wire  regs_234_clock;
  wire  regs_234_reset;
  wire [63:0] regs_234_io_in;
  wire [63:0] regs_234_io_init;
  wire  regs_234_io_reset;
  wire [63:0] regs_234_io_out;
  wire  regs_234_io_enable;
  wire  regs_235_clock;
  wire  regs_235_reset;
  wire [63:0] regs_235_io_in;
  wire [63:0] regs_235_io_init;
  wire  regs_235_io_reset;
  wire [63:0] regs_235_io_out;
  wire  regs_235_io_enable;
  wire  regs_236_clock;
  wire  regs_236_reset;
  wire [63:0] regs_236_io_in;
  wire [63:0] regs_236_io_init;
  wire  regs_236_io_reset;
  wire [63:0] regs_236_io_out;
  wire  regs_236_io_enable;
  wire  regs_237_clock;
  wire  regs_237_reset;
  wire [63:0] regs_237_io_in;
  wire [63:0] regs_237_io_init;
  wire  regs_237_io_reset;
  wire [63:0] regs_237_io_out;
  wire  regs_237_io_enable;
  wire  regs_238_clock;
  wire  regs_238_reset;
  wire [63:0] regs_238_io_in;
  wire [63:0] regs_238_io_init;
  wire  regs_238_io_reset;
  wire [63:0] regs_238_io_out;
  wire  regs_238_io_enable;
  wire  regs_239_clock;
  wire  regs_239_reset;
  wire [63:0] regs_239_io_in;
  wire [63:0] regs_239_io_init;
  wire  regs_239_io_reset;
  wire [63:0] regs_239_io_out;
  wire  regs_239_io_enable;
  wire  regs_240_clock;
  wire  regs_240_reset;
  wire [63:0] regs_240_io_in;
  wire [63:0] regs_240_io_init;
  wire  regs_240_io_reset;
  wire [63:0] regs_240_io_out;
  wire  regs_240_io_enable;
  wire  regs_241_clock;
  wire  regs_241_reset;
  wire [63:0] regs_241_io_in;
  wire [63:0] regs_241_io_init;
  wire  regs_241_io_reset;
  wire [63:0] regs_241_io_out;
  wire  regs_241_io_enable;
  wire  regs_242_clock;
  wire  regs_242_reset;
  wire [63:0] regs_242_io_in;
  wire [63:0] regs_242_io_init;
  wire  regs_242_io_reset;
  wire [63:0] regs_242_io_out;
  wire  regs_242_io_enable;
  wire  regs_243_clock;
  wire  regs_243_reset;
  wire [63:0] regs_243_io_in;
  wire [63:0] regs_243_io_init;
  wire  regs_243_io_reset;
  wire [63:0] regs_243_io_out;
  wire  regs_243_io_enable;
  wire  regs_244_clock;
  wire  regs_244_reset;
  wire [63:0] regs_244_io_in;
  wire [63:0] regs_244_io_init;
  wire  regs_244_io_reset;
  wire [63:0] regs_244_io_out;
  wire  regs_244_io_enable;
  wire  regs_245_clock;
  wire  regs_245_reset;
  wire [63:0] regs_245_io_in;
  wire [63:0] regs_245_io_init;
  wire  regs_245_io_reset;
  wire [63:0] regs_245_io_out;
  wire  regs_245_io_enable;
  wire  regs_246_clock;
  wire  regs_246_reset;
  wire [63:0] regs_246_io_in;
  wire [63:0] regs_246_io_init;
  wire  regs_246_io_reset;
  wire [63:0] regs_246_io_out;
  wire  regs_246_io_enable;
  wire  regs_247_clock;
  wire  regs_247_reset;
  wire [63:0] regs_247_io_in;
  wire [63:0] regs_247_io_init;
  wire  regs_247_io_reset;
  wire [63:0] regs_247_io_out;
  wire  regs_247_io_enable;
  wire  regs_248_clock;
  wire  regs_248_reset;
  wire [63:0] regs_248_io_in;
  wire [63:0] regs_248_io_init;
  wire  regs_248_io_reset;
  wire [63:0] regs_248_io_out;
  wire  regs_248_io_enable;
  wire  regs_249_clock;
  wire  regs_249_reset;
  wire [63:0] regs_249_io_in;
  wire [63:0] regs_249_io_init;
  wire  regs_249_io_reset;
  wire [63:0] regs_249_io_out;
  wire  regs_249_io_enable;
  wire  regs_250_clock;
  wire  regs_250_reset;
  wire [63:0] regs_250_io_in;
  wire [63:0] regs_250_io_init;
  wire  regs_250_io_reset;
  wire [63:0] regs_250_io_out;
  wire  regs_250_io_enable;
  wire  regs_251_clock;
  wire  regs_251_reset;
  wire [63:0] regs_251_io_in;
  wire [63:0] regs_251_io_init;
  wire  regs_251_io_reset;
  wire [63:0] regs_251_io_out;
  wire  regs_251_io_enable;
  wire  regs_252_clock;
  wire  regs_252_reset;
  wire [63:0] regs_252_io_in;
  wire [63:0] regs_252_io_init;
  wire  regs_252_io_reset;
  wire [63:0] regs_252_io_out;
  wire  regs_252_io_enable;
  wire  regs_253_clock;
  wire  regs_253_reset;
  wire [63:0] regs_253_io_in;
  wire [63:0] regs_253_io_init;
  wire  regs_253_io_reset;
  wire [63:0] regs_253_io_out;
  wire  regs_253_io_enable;
  wire  regs_254_clock;
  wire  regs_254_reset;
  wire [63:0] regs_254_io_in;
  wire [63:0] regs_254_io_init;
  wire  regs_254_io_reset;
  wire [63:0] regs_254_io_out;
  wire  regs_254_io_enable;
  wire  regs_255_clock;
  wire  regs_255_reset;
  wire [63:0] regs_255_io_in;
  wire [63:0] regs_255_io_init;
  wire  regs_255_io_reset;
  wire [63:0] regs_255_io_out;
  wire  regs_255_io_enable;
  wire  regs_256_clock;
  wire  regs_256_reset;
  wire [63:0] regs_256_io_in;
  wire [63:0] regs_256_io_init;
  wire  regs_256_io_reset;
  wire [63:0] regs_256_io_out;
  wire  regs_256_io_enable;
  wire  regs_257_clock;
  wire  regs_257_reset;
  wire [63:0] regs_257_io_in;
  wire [63:0] regs_257_io_init;
  wire  regs_257_io_reset;
  wire [63:0] regs_257_io_out;
  wire  regs_257_io_enable;
  wire  regs_258_clock;
  wire  regs_258_reset;
  wire [63:0] regs_258_io_in;
  wire [63:0] regs_258_io_init;
  wire  regs_258_io_reset;
  wire [63:0] regs_258_io_out;
  wire  regs_258_io_enable;
  wire  regs_259_clock;
  wire  regs_259_reset;
  wire [63:0] regs_259_io_in;
  wire [63:0] regs_259_io_init;
  wire  regs_259_io_reset;
  wire [63:0] regs_259_io_out;
  wire  regs_259_io_enable;
  wire  regs_260_clock;
  wire  regs_260_reset;
  wire [63:0] regs_260_io_in;
  wire [63:0] regs_260_io_init;
  wire  regs_260_io_reset;
  wire [63:0] regs_260_io_out;
  wire  regs_260_io_enable;
  wire  regs_261_clock;
  wire  regs_261_reset;
  wire [63:0] regs_261_io_in;
  wire [63:0] regs_261_io_init;
  wire  regs_261_io_reset;
  wire [63:0] regs_261_io_out;
  wire  regs_261_io_enable;
  wire  regs_262_clock;
  wire  regs_262_reset;
  wire [63:0] regs_262_io_in;
  wire [63:0] regs_262_io_init;
  wire  regs_262_io_reset;
  wire [63:0] regs_262_io_out;
  wire  regs_262_io_enable;
  wire  regs_263_clock;
  wire  regs_263_reset;
  wire [63:0] regs_263_io_in;
  wire [63:0] regs_263_io_init;
  wire  regs_263_io_reset;
  wire [63:0] regs_263_io_out;
  wire  regs_263_io_enable;
  wire  regs_264_clock;
  wire  regs_264_reset;
  wire [63:0] regs_264_io_in;
  wire [63:0] regs_264_io_init;
  wire  regs_264_io_reset;
  wire [63:0] regs_264_io_out;
  wire  regs_264_io_enable;
  wire  regs_265_clock;
  wire  regs_265_reset;
  wire [63:0] regs_265_io_in;
  wire [63:0] regs_265_io_init;
  wire  regs_265_io_reset;
  wire [63:0] regs_265_io_out;
  wire  regs_265_io_enable;
  wire  regs_266_clock;
  wire  regs_266_reset;
  wire [63:0] regs_266_io_in;
  wire [63:0] regs_266_io_init;
  wire  regs_266_io_reset;
  wire [63:0] regs_266_io_out;
  wire  regs_266_io_enable;
  wire  regs_267_clock;
  wire  regs_267_reset;
  wire [63:0] regs_267_io_in;
  wire [63:0] regs_267_io_init;
  wire  regs_267_io_reset;
  wire [63:0] regs_267_io_out;
  wire  regs_267_io_enable;
  wire  regs_268_clock;
  wire  regs_268_reset;
  wire [63:0] regs_268_io_in;
  wire [63:0] regs_268_io_init;
  wire  regs_268_io_reset;
  wire [63:0] regs_268_io_out;
  wire  regs_268_io_enable;
  wire  regs_269_clock;
  wire  regs_269_reset;
  wire [63:0] regs_269_io_in;
  wire [63:0] regs_269_io_init;
  wire  regs_269_io_reset;
  wire [63:0] regs_269_io_out;
  wire  regs_269_io_enable;
  wire  regs_270_clock;
  wire  regs_270_reset;
  wire [63:0] regs_270_io_in;
  wire [63:0] regs_270_io_init;
  wire  regs_270_io_reset;
  wire [63:0] regs_270_io_out;
  wire  regs_270_io_enable;
  wire  regs_271_clock;
  wire  regs_271_reset;
  wire [63:0] regs_271_io_in;
  wire [63:0] regs_271_io_init;
  wire  regs_271_io_reset;
  wire [63:0] regs_271_io_out;
  wire  regs_271_io_enable;
  wire  regs_272_clock;
  wire  regs_272_reset;
  wire [63:0] regs_272_io_in;
  wire [63:0] regs_272_io_init;
  wire  regs_272_io_reset;
  wire [63:0] regs_272_io_out;
  wire  regs_272_io_enable;
  wire  regs_273_clock;
  wire  regs_273_reset;
  wire [63:0] regs_273_io_in;
  wire [63:0] regs_273_io_init;
  wire  regs_273_io_reset;
  wire [63:0] regs_273_io_out;
  wire  regs_273_io_enable;
  wire  regs_274_clock;
  wire  regs_274_reset;
  wire [63:0] regs_274_io_in;
  wire [63:0] regs_274_io_init;
  wire  regs_274_io_reset;
  wire [63:0] regs_274_io_out;
  wire  regs_274_io_enable;
  wire  regs_275_clock;
  wire  regs_275_reset;
  wire [63:0] regs_275_io_in;
  wire [63:0] regs_275_io_init;
  wire  regs_275_io_reset;
  wire [63:0] regs_275_io_out;
  wire  regs_275_io_enable;
  wire  regs_276_clock;
  wire  regs_276_reset;
  wire [63:0] regs_276_io_in;
  wire [63:0] regs_276_io_init;
  wire  regs_276_io_reset;
  wire [63:0] regs_276_io_out;
  wire  regs_276_io_enable;
  wire  regs_277_clock;
  wire  regs_277_reset;
  wire [63:0] regs_277_io_in;
  wire [63:0] regs_277_io_init;
  wire  regs_277_io_reset;
  wire [63:0] regs_277_io_out;
  wire  regs_277_io_enable;
  wire  regs_278_clock;
  wire  regs_278_reset;
  wire [63:0] regs_278_io_in;
  wire [63:0] regs_278_io_init;
  wire  regs_278_io_reset;
  wire [63:0] regs_278_io_out;
  wire  regs_278_io_enable;
  wire  regs_279_clock;
  wire  regs_279_reset;
  wire [63:0] regs_279_io_in;
  wire [63:0] regs_279_io_init;
  wire  regs_279_io_reset;
  wire [63:0] regs_279_io_out;
  wire  regs_279_io_enable;
  wire  regs_280_clock;
  wire  regs_280_reset;
  wire [63:0] regs_280_io_in;
  wire [63:0] regs_280_io_init;
  wire  regs_280_io_reset;
  wire [63:0] regs_280_io_out;
  wire  regs_280_io_enable;
  wire  regs_281_clock;
  wire  regs_281_reset;
  wire [63:0] regs_281_io_in;
  wire [63:0] regs_281_io_init;
  wire  regs_281_io_reset;
  wire [63:0] regs_281_io_out;
  wire  regs_281_io_enable;
  wire  regs_282_clock;
  wire  regs_282_reset;
  wire [63:0] regs_282_io_in;
  wire [63:0] regs_282_io_init;
  wire  regs_282_io_reset;
  wire [63:0] regs_282_io_out;
  wire  regs_282_io_enable;
  wire  regs_283_clock;
  wire  regs_283_reset;
  wire [63:0] regs_283_io_in;
  wire [63:0] regs_283_io_init;
  wire  regs_283_io_reset;
  wire [63:0] regs_283_io_out;
  wire  regs_283_io_enable;
  wire  regs_284_clock;
  wire  regs_284_reset;
  wire [63:0] regs_284_io_in;
  wire [63:0] regs_284_io_init;
  wire  regs_284_io_reset;
  wire [63:0] regs_284_io_out;
  wire  regs_284_io_enable;
  wire  regs_285_clock;
  wire  regs_285_reset;
  wire [63:0] regs_285_io_in;
  wire [63:0] regs_285_io_init;
  wire  regs_285_io_reset;
  wire [63:0] regs_285_io_out;
  wire  regs_285_io_enable;
  wire  regs_286_clock;
  wire  regs_286_reset;
  wire [63:0] regs_286_io_in;
  wire [63:0] regs_286_io_init;
  wire  regs_286_io_reset;
  wire [63:0] regs_286_io_out;
  wire  regs_286_io_enable;
  wire  regs_287_clock;
  wire  regs_287_reset;
  wire [63:0] regs_287_io_in;
  wire [63:0] regs_287_io_init;
  wire  regs_287_io_reset;
  wire [63:0] regs_287_io_out;
  wire  regs_287_io_enable;
  wire  regs_288_clock;
  wire  regs_288_reset;
  wire [63:0] regs_288_io_in;
  wire [63:0] regs_288_io_init;
  wire  regs_288_io_reset;
  wire [63:0] regs_288_io_out;
  wire  regs_288_io_enable;
  wire  regs_289_clock;
  wire  regs_289_reset;
  wire [63:0] regs_289_io_in;
  wire [63:0] regs_289_io_init;
  wire  regs_289_io_reset;
  wire [63:0] regs_289_io_out;
  wire  regs_289_io_enable;
  wire  regs_290_clock;
  wire  regs_290_reset;
  wire [63:0] regs_290_io_in;
  wire [63:0] regs_290_io_init;
  wire  regs_290_io_reset;
  wire [63:0] regs_290_io_out;
  wire  regs_290_io_enable;
  wire  regs_291_clock;
  wire  regs_291_reset;
  wire [63:0] regs_291_io_in;
  wire [63:0] regs_291_io_init;
  wire  regs_291_io_reset;
  wire [63:0] regs_291_io_out;
  wire  regs_291_io_enable;
  wire  regs_292_clock;
  wire  regs_292_reset;
  wire [63:0] regs_292_io_in;
  wire [63:0] regs_292_io_init;
  wire  regs_292_io_reset;
  wire [63:0] regs_292_io_out;
  wire  regs_292_io_enable;
  wire  regs_293_clock;
  wire  regs_293_reset;
  wire [63:0] regs_293_io_in;
  wire [63:0] regs_293_io_init;
  wire  regs_293_io_reset;
  wire [63:0] regs_293_io_out;
  wire  regs_293_io_enable;
  wire  regs_294_clock;
  wire  regs_294_reset;
  wire [63:0] regs_294_io_in;
  wire [63:0] regs_294_io_init;
  wire  regs_294_io_reset;
  wire [63:0] regs_294_io_out;
  wire  regs_294_io_enable;
  wire  regs_295_clock;
  wire  regs_295_reset;
  wire [63:0] regs_295_io_in;
  wire [63:0] regs_295_io_init;
  wire  regs_295_io_reset;
  wire [63:0] regs_295_io_out;
  wire  regs_295_io_enable;
  wire  regs_296_clock;
  wire  regs_296_reset;
  wire [63:0] regs_296_io_in;
  wire [63:0] regs_296_io_init;
  wire  regs_296_io_reset;
  wire [63:0] regs_296_io_out;
  wire  regs_296_io_enable;
  wire  regs_297_clock;
  wire  regs_297_reset;
  wire [63:0] regs_297_io_in;
  wire [63:0] regs_297_io_init;
  wire  regs_297_io_reset;
  wire [63:0] regs_297_io_out;
  wire  regs_297_io_enable;
  wire  regs_298_clock;
  wire  regs_298_reset;
  wire [63:0] regs_298_io_in;
  wire [63:0] regs_298_io_init;
  wire  regs_298_io_reset;
  wire [63:0] regs_298_io_out;
  wire  regs_298_io_enable;
  wire  regs_299_clock;
  wire  regs_299_reset;
  wire [63:0] regs_299_io_in;
  wire [63:0] regs_299_io_init;
  wire  regs_299_io_reset;
  wire [63:0] regs_299_io_out;
  wire  regs_299_io_enable;
  wire  regs_300_clock;
  wire  regs_300_reset;
  wire [63:0] regs_300_io_in;
  wire [63:0] regs_300_io_init;
  wire  regs_300_io_reset;
  wire [63:0] regs_300_io_out;
  wire  regs_300_io_enable;
  wire  regs_301_clock;
  wire  regs_301_reset;
  wire [63:0] regs_301_io_in;
  wire [63:0] regs_301_io_init;
  wire  regs_301_io_reset;
  wire [63:0] regs_301_io_out;
  wire  regs_301_io_enable;
  wire  regs_302_clock;
  wire  regs_302_reset;
  wire [63:0] regs_302_io_in;
  wire [63:0] regs_302_io_init;
  wire  regs_302_io_reset;
  wire [63:0] regs_302_io_out;
  wire  regs_302_io_enable;
  wire  regs_303_clock;
  wire  regs_303_reset;
  wire [63:0] regs_303_io_in;
  wire [63:0] regs_303_io_init;
  wire  regs_303_io_reset;
  wire [63:0] regs_303_io_out;
  wire  regs_303_io_enable;
  wire  regs_304_clock;
  wire  regs_304_reset;
  wire [63:0] regs_304_io_in;
  wire [63:0] regs_304_io_init;
  wire  regs_304_io_reset;
  wire [63:0] regs_304_io_out;
  wire  regs_304_io_enable;
  wire  regs_305_clock;
  wire  regs_305_reset;
  wire [63:0] regs_305_io_in;
  wire [63:0] regs_305_io_init;
  wire  regs_305_io_reset;
  wire [63:0] regs_305_io_out;
  wire  regs_305_io_enable;
  wire  regs_306_clock;
  wire  regs_306_reset;
  wire [63:0] regs_306_io_in;
  wire [63:0] regs_306_io_init;
  wire  regs_306_io_reset;
  wire [63:0] regs_306_io_out;
  wire  regs_306_io_enable;
  wire  regs_307_clock;
  wire  regs_307_reset;
  wire [63:0] regs_307_io_in;
  wire [63:0] regs_307_io_init;
  wire  regs_307_io_reset;
  wire [63:0] regs_307_io_out;
  wire  regs_307_io_enable;
  wire  regs_308_clock;
  wire  regs_308_reset;
  wire [63:0] regs_308_io_in;
  wire [63:0] regs_308_io_init;
  wire  regs_308_io_reset;
  wire [63:0] regs_308_io_out;
  wire  regs_308_io_enable;
  wire  regs_309_clock;
  wire  regs_309_reset;
  wire [63:0] regs_309_io_in;
  wire [63:0] regs_309_io_init;
  wire  regs_309_io_reset;
  wire [63:0] regs_309_io_out;
  wire  regs_309_io_enable;
  wire  regs_310_clock;
  wire  regs_310_reset;
  wire [63:0] regs_310_io_in;
  wire [63:0] regs_310_io_init;
  wire  regs_310_io_reset;
  wire [63:0] regs_310_io_out;
  wire  regs_310_io_enable;
  wire  regs_311_clock;
  wire  regs_311_reset;
  wire [63:0] regs_311_io_in;
  wire [63:0] regs_311_io_init;
  wire  regs_311_io_reset;
  wire [63:0] regs_311_io_out;
  wire  regs_311_io_enable;
  wire  regs_312_clock;
  wire  regs_312_reset;
  wire [63:0] regs_312_io_in;
  wire [63:0] regs_312_io_init;
  wire  regs_312_io_reset;
  wire [63:0] regs_312_io_out;
  wire  regs_312_io_enable;
  wire  regs_313_clock;
  wire  regs_313_reset;
  wire [63:0] regs_313_io_in;
  wire [63:0] regs_313_io_init;
  wire  regs_313_io_reset;
  wire [63:0] regs_313_io_out;
  wire  regs_313_io_enable;
  wire  regs_314_clock;
  wire  regs_314_reset;
  wire [63:0] regs_314_io_in;
  wire [63:0] regs_314_io_init;
  wire  regs_314_io_reset;
  wire [63:0] regs_314_io_out;
  wire  regs_314_io_enable;
  wire  regs_315_clock;
  wire  regs_315_reset;
  wire [63:0] regs_315_io_in;
  wire [63:0] regs_315_io_init;
  wire  regs_315_io_reset;
  wire [63:0] regs_315_io_out;
  wire  regs_315_io_enable;
  wire  regs_316_clock;
  wire  regs_316_reset;
  wire [63:0] regs_316_io_in;
  wire [63:0] regs_316_io_init;
  wire  regs_316_io_reset;
  wire [63:0] regs_316_io_out;
  wire  regs_316_io_enable;
  wire  regs_317_clock;
  wire  regs_317_reset;
  wire [63:0] regs_317_io_in;
  wire [63:0] regs_317_io_init;
  wire  regs_317_io_reset;
  wire [63:0] regs_317_io_out;
  wire  regs_317_io_enable;
  wire  regs_318_clock;
  wire  regs_318_reset;
  wire [63:0] regs_318_io_in;
  wire [63:0] regs_318_io_init;
  wire  regs_318_io_reset;
  wire [63:0] regs_318_io_out;
  wire  regs_318_io_enable;
  wire  regs_319_clock;
  wire  regs_319_reset;
  wire [63:0] regs_319_io_in;
  wire [63:0] regs_319_io_init;
  wire  regs_319_io_reset;
  wire [63:0] regs_319_io_out;
  wire  regs_319_io_enable;
  wire  regs_320_clock;
  wire  regs_320_reset;
  wire [63:0] regs_320_io_in;
  wire [63:0] regs_320_io_init;
  wire  regs_320_io_reset;
  wire [63:0] regs_320_io_out;
  wire  regs_320_io_enable;
  wire  regs_321_clock;
  wire  regs_321_reset;
  wire [63:0] regs_321_io_in;
  wire [63:0] regs_321_io_init;
  wire  regs_321_io_reset;
  wire [63:0] regs_321_io_out;
  wire  regs_321_io_enable;
  wire  regs_322_clock;
  wire  regs_322_reset;
  wire [63:0] regs_322_io_in;
  wire [63:0] regs_322_io_init;
  wire  regs_322_io_reset;
  wire [63:0] regs_322_io_out;
  wire  regs_322_io_enable;
  wire  regs_323_clock;
  wire  regs_323_reset;
  wire [63:0] regs_323_io_in;
  wire [63:0] regs_323_io_init;
  wire  regs_323_io_reset;
  wire [63:0] regs_323_io_out;
  wire  regs_323_io_enable;
  wire  regs_324_clock;
  wire  regs_324_reset;
  wire [63:0] regs_324_io_in;
  wire [63:0] regs_324_io_init;
  wire  regs_324_io_reset;
  wire [63:0] regs_324_io_out;
  wire  regs_324_io_enable;
  wire  regs_325_clock;
  wire  regs_325_reset;
  wire [63:0] regs_325_io_in;
  wire [63:0] regs_325_io_init;
  wire  regs_325_io_reset;
  wire [63:0] regs_325_io_out;
  wire  regs_325_io_enable;
  wire  regs_326_clock;
  wire  regs_326_reset;
  wire [63:0] regs_326_io_in;
  wire [63:0] regs_326_io_init;
  wire  regs_326_io_reset;
  wire [63:0] regs_326_io_out;
  wire  regs_326_io_enable;
  wire  regs_327_clock;
  wire  regs_327_reset;
  wire [63:0] regs_327_io_in;
  wire [63:0] regs_327_io_init;
  wire  regs_327_io_reset;
  wire [63:0] regs_327_io_out;
  wire  regs_327_io_enable;
  wire  regs_328_clock;
  wire  regs_328_reset;
  wire [63:0] regs_328_io_in;
  wire [63:0] regs_328_io_init;
  wire  regs_328_io_reset;
  wire [63:0] regs_328_io_out;
  wire  regs_328_io_enable;
  wire  regs_329_clock;
  wire  regs_329_reset;
  wire [63:0] regs_329_io_in;
  wire [63:0] regs_329_io_init;
  wire  regs_329_io_reset;
  wire [63:0] regs_329_io_out;
  wire  regs_329_io_enable;
  wire  regs_330_clock;
  wire  regs_330_reset;
  wire [63:0] regs_330_io_in;
  wire [63:0] regs_330_io_init;
  wire  regs_330_io_reset;
  wire [63:0] regs_330_io_out;
  wire  regs_330_io_enable;
  wire  regs_331_clock;
  wire  regs_331_reset;
  wire [63:0] regs_331_io_in;
  wire [63:0] regs_331_io_init;
  wire  regs_331_io_reset;
  wire [63:0] regs_331_io_out;
  wire  regs_331_io_enable;
  wire  regs_332_clock;
  wire  regs_332_reset;
  wire [63:0] regs_332_io_in;
  wire [63:0] regs_332_io_init;
  wire  regs_332_io_reset;
  wire [63:0] regs_332_io_out;
  wire  regs_332_io_enable;
  wire  regs_333_clock;
  wire  regs_333_reset;
  wire [63:0] regs_333_io_in;
  wire [63:0] regs_333_io_init;
  wire  regs_333_io_reset;
  wire [63:0] regs_333_io_out;
  wire  regs_333_io_enable;
  wire  regs_334_clock;
  wire  regs_334_reset;
  wire [63:0] regs_334_io_in;
  wire [63:0] regs_334_io_init;
  wire  regs_334_io_reset;
  wire [63:0] regs_334_io_out;
  wire  regs_334_io_enable;
  wire  regs_335_clock;
  wire  regs_335_reset;
  wire [63:0] regs_335_io_in;
  wire [63:0] regs_335_io_init;
  wire  regs_335_io_reset;
  wire [63:0] regs_335_io_out;
  wire  regs_335_io_enable;
  wire  regs_336_clock;
  wire  regs_336_reset;
  wire [63:0] regs_336_io_in;
  wire [63:0] regs_336_io_init;
  wire  regs_336_io_reset;
  wire [63:0] regs_336_io_out;
  wire  regs_336_io_enable;
  wire  regs_337_clock;
  wire  regs_337_reset;
  wire [63:0] regs_337_io_in;
  wire [63:0] regs_337_io_init;
  wire  regs_337_io_reset;
  wire [63:0] regs_337_io_out;
  wire  regs_337_io_enable;
  wire  regs_338_clock;
  wire  regs_338_reset;
  wire [63:0] regs_338_io_in;
  wire [63:0] regs_338_io_init;
  wire  regs_338_io_reset;
  wire [63:0] regs_338_io_out;
  wire  regs_338_io_enable;
  wire  regs_339_clock;
  wire  regs_339_reset;
  wire [63:0] regs_339_io_in;
  wire [63:0] regs_339_io_init;
  wire  regs_339_io_reset;
  wire [63:0] regs_339_io_out;
  wire  regs_339_io_enable;
  wire  regs_340_clock;
  wire  regs_340_reset;
  wire [63:0] regs_340_io_in;
  wire [63:0] regs_340_io_init;
  wire  regs_340_io_reset;
  wire [63:0] regs_340_io_out;
  wire  regs_340_io_enable;
  wire  regs_341_clock;
  wire  regs_341_reset;
  wire [63:0] regs_341_io_in;
  wire [63:0] regs_341_io_init;
  wire  regs_341_io_reset;
  wire [63:0] regs_341_io_out;
  wire  regs_341_io_enable;
  wire  regs_342_clock;
  wire  regs_342_reset;
  wire [63:0] regs_342_io_in;
  wire [63:0] regs_342_io_init;
  wire  regs_342_io_reset;
  wire [63:0] regs_342_io_out;
  wire  regs_342_io_enable;
  wire  regs_343_clock;
  wire  regs_343_reset;
  wire [63:0] regs_343_io_in;
  wire [63:0] regs_343_io_init;
  wire  regs_343_io_reset;
  wire [63:0] regs_343_io_out;
  wire  regs_343_io_enable;
  wire  regs_344_clock;
  wire  regs_344_reset;
  wire [63:0] regs_344_io_in;
  wire [63:0] regs_344_io_init;
  wire  regs_344_io_reset;
  wire [63:0] regs_344_io_out;
  wire  regs_344_io_enable;
  wire  regs_345_clock;
  wire  regs_345_reset;
  wire [63:0] regs_345_io_in;
  wire [63:0] regs_345_io_init;
  wire  regs_345_io_reset;
  wire [63:0] regs_345_io_out;
  wire  regs_345_io_enable;
  wire  regs_346_clock;
  wire  regs_346_reset;
  wire [63:0] regs_346_io_in;
  wire [63:0] regs_346_io_init;
  wire  regs_346_io_reset;
  wire [63:0] regs_346_io_out;
  wire  regs_346_io_enable;
  wire  regs_347_clock;
  wire  regs_347_reset;
  wire [63:0] regs_347_io_in;
  wire [63:0] regs_347_io_init;
  wire  regs_347_io_reset;
  wire [63:0] regs_347_io_out;
  wire  regs_347_io_enable;
  wire  regs_348_clock;
  wire  regs_348_reset;
  wire [63:0] regs_348_io_in;
  wire [63:0] regs_348_io_init;
  wire  regs_348_io_reset;
  wire [63:0] regs_348_io_out;
  wire  regs_348_io_enable;
  wire  regs_349_clock;
  wire  regs_349_reset;
  wire [63:0] regs_349_io_in;
  wire [63:0] regs_349_io_init;
  wire  regs_349_io_reset;
  wire [63:0] regs_349_io_out;
  wire  regs_349_io_enable;
  wire  regs_350_clock;
  wire  regs_350_reset;
  wire [63:0] regs_350_io_in;
  wire [63:0] regs_350_io_init;
  wire  regs_350_io_reset;
  wire [63:0] regs_350_io_out;
  wire  regs_350_io_enable;
  wire  regs_351_clock;
  wire  regs_351_reset;
  wire [63:0] regs_351_io_in;
  wire [63:0] regs_351_io_init;
  wire  regs_351_io_reset;
  wire [63:0] regs_351_io_out;
  wire  regs_351_io_enable;
  wire  regs_352_clock;
  wire  regs_352_reset;
  wire [63:0] regs_352_io_in;
  wire [63:0] regs_352_io_init;
  wire  regs_352_io_reset;
  wire [63:0] regs_352_io_out;
  wire  regs_352_io_enable;
  wire  regs_353_clock;
  wire  regs_353_reset;
  wire [63:0] regs_353_io_in;
  wire [63:0] regs_353_io_init;
  wire  regs_353_io_reset;
  wire [63:0] regs_353_io_out;
  wire  regs_353_io_enable;
  wire  regs_354_clock;
  wire  regs_354_reset;
  wire [63:0] regs_354_io_in;
  wire [63:0] regs_354_io_init;
  wire  regs_354_io_reset;
  wire [63:0] regs_354_io_out;
  wire  regs_354_io_enable;
  wire  regs_355_clock;
  wire  regs_355_reset;
  wire [63:0] regs_355_io_in;
  wire [63:0] regs_355_io_init;
  wire  regs_355_io_reset;
  wire [63:0] regs_355_io_out;
  wire  regs_355_io_enable;
  wire  regs_356_clock;
  wire  regs_356_reset;
  wire [63:0] regs_356_io_in;
  wire [63:0] regs_356_io_init;
  wire  regs_356_io_reset;
  wire [63:0] regs_356_io_out;
  wire  regs_356_io_enable;
  wire  regs_357_clock;
  wire  regs_357_reset;
  wire [63:0] regs_357_io_in;
  wire [63:0] regs_357_io_init;
  wire  regs_357_io_reset;
  wire [63:0] regs_357_io_out;
  wire  regs_357_io_enable;
  wire  regs_358_clock;
  wire  regs_358_reset;
  wire [63:0] regs_358_io_in;
  wire [63:0] regs_358_io_init;
  wire  regs_358_io_reset;
  wire [63:0] regs_358_io_out;
  wire  regs_358_io_enable;
  wire  regs_359_clock;
  wire  regs_359_reset;
  wire [63:0] regs_359_io_in;
  wire [63:0] regs_359_io_init;
  wire  regs_359_io_reset;
  wire [63:0] regs_359_io_out;
  wire  regs_359_io_enable;
  wire  regs_360_clock;
  wire  regs_360_reset;
  wire [63:0] regs_360_io_in;
  wire [63:0] regs_360_io_init;
  wire  regs_360_io_reset;
  wire [63:0] regs_360_io_out;
  wire  regs_360_io_enable;
  wire  regs_361_clock;
  wire  regs_361_reset;
  wire [63:0] regs_361_io_in;
  wire [63:0] regs_361_io_init;
  wire  regs_361_io_reset;
  wire [63:0] regs_361_io_out;
  wire  regs_361_io_enable;
  wire  regs_362_clock;
  wire  regs_362_reset;
  wire [63:0] regs_362_io_in;
  wire [63:0] regs_362_io_init;
  wire  regs_362_io_reset;
  wire [63:0] regs_362_io_out;
  wire  regs_362_io_enable;
  wire  regs_363_clock;
  wire  regs_363_reset;
  wire [63:0] regs_363_io_in;
  wire [63:0] regs_363_io_init;
  wire  regs_363_io_reset;
  wire [63:0] regs_363_io_out;
  wire  regs_363_io_enable;
  wire  regs_364_clock;
  wire  regs_364_reset;
  wire [63:0] regs_364_io_in;
  wire [63:0] regs_364_io_init;
  wire  regs_364_io_reset;
  wire [63:0] regs_364_io_out;
  wire  regs_364_io_enable;
  wire  regs_365_clock;
  wire  regs_365_reset;
  wire [63:0] regs_365_io_in;
  wire [63:0] regs_365_io_init;
  wire  regs_365_io_reset;
  wire [63:0] regs_365_io_out;
  wire  regs_365_io_enable;
  wire  regs_366_clock;
  wire  regs_366_reset;
  wire [63:0] regs_366_io_in;
  wire [63:0] regs_366_io_init;
  wire  regs_366_io_reset;
  wire [63:0] regs_366_io_out;
  wire  regs_366_io_enable;
  wire  regs_367_clock;
  wire  regs_367_reset;
  wire [63:0] regs_367_io_in;
  wire [63:0] regs_367_io_init;
  wire  regs_367_io_reset;
  wire [63:0] regs_367_io_out;
  wire  regs_367_io_enable;
  wire  regs_368_clock;
  wire  regs_368_reset;
  wire [63:0] regs_368_io_in;
  wire [63:0] regs_368_io_init;
  wire  regs_368_io_reset;
  wire [63:0] regs_368_io_out;
  wire  regs_368_io_enable;
  wire  regs_369_clock;
  wire  regs_369_reset;
  wire [63:0] regs_369_io_in;
  wire [63:0] regs_369_io_init;
  wire  regs_369_io_reset;
  wire [63:0] regs_369_io_out;
  wire  regs_369_io_enable;
  wire  regs_370_clock;
  wire  regs_370_reset;
  wire [63:0] regs_370_io_in;
  wire [63:0] regs_370_io_init;
  wire  regs_370_io_reset;
  wire [63:0] regs_370_io_out;
  wire  regs_370_io_enable;
  wire  regs_371_clock;
  wire  regs_371_reset;
  wire [63:0] regs_371_io_in;
  wire [63:0] regs_371_io_init;
  wire  regs_371_io_reset;
  wire [63:0] regs_371_io_out;
  wire  regs_371_io_enable;
  wire  regs_372_clock;
  wire  regs_372_reset;
  wire [63:0] regs_372_io_in;
  wire [63:0] regs_372_io_init;
  wire  regs_372_io_reset;
  wire [63:0] regs_372_io_out;
  wire  regs_372_io_enable;
  wire  regs_373_clock;
  wire  regs_373_reset;
  wire [63:0] regs_373_io_in;
  wire [63:0] regs_373_io_init;
  wire  regs_373_io_reset;
  wire [63:0] regs_373_io_out;
  wire  regs_373_io_enable;
  wire  regs_374_clock;
  wire  regs_374_reset;
  wire [63:0] regs_374_io_in;
  wire [63:0] regs_374_io_init;
  wire  regs_374_io_reset;
  wire [63:0] regs_374_io_out;
  wire  regs_374_io_enable;
  wire  regs_375_clock;
  wire  regs_375_reset;
  wire [63:0] regs_375_io_in;
  wire [63:0] regs_375_io_init;
  wire  regs_375_io_reset;
  wire [63:0] regs_375_io_out;
  wire  regs_375_io_enable;
  wire  regs_376_clock;
  wire  regs_376_reset;
  wire [63:0] regs_376_io_in;
  wire [63:0] regs_376_io_init;
  wire  regs_376_io_reset;
  wire [63:0] regs_376_io_out;
  wire  regs_376_io_enable;
  wire  regs_377_clock;
  wire  regs_377_reset;
  wire [63:0] regs_377_io_in;
  wire [63:0] regs_377_io_init;
  wire  regs_377_io_reset;
  wire [63:0] regs_377_io_out;
  wire  regs_377_io_enable;
  wire  regs_378_clock;
  wire  regs_378_reset;
  wire [63:0] regs_378_io_in;
  wire [63:0] regs_378_io_init;
  wire  regs_378_io_reset;
  wire [63:0] regs_378_io_out;
  wire  regs_378_io_enable;
  wire  regs_379_clock;
  wire  regs_379_reset;
  wire [63:0] regs_379_io_in;
  wire [63:0] regs_379_io_init;
  wire  regs_379_io_reset;
  wire [63:0] regs_379_io_out;
  wire  regs_379_io_enable;
  wire  regs_380_clock;
  wire  regs_380_reset;
  wire [63:0] regs_380_io_in;
  wire [63:0] regs_380_io_init;
  wire  regs_380_io_reset;
  wire [63:0] regs_380_io_out;
  wire  regs_380_io_enable;
  wire  regs_381_clock;
  wire  regs_381_reset;
  wire [63:0] regs_381_io_in;
  wire [63:0] regs_381_io_init;
  wire  regs_381_io_reset;
  wire [63:0] regs_381_io_out;
  wire  regs_381_io_enable;
  wire  regs_382_clock;
  wire  regs_382_reset;
  wire [63:0] regs_382_io_in;
  wire [63:0] regs_382_io_init;
  wire  regs_382_io_reset;
  wire [63:0] regs_382_io_out;
  wire  regs_382_io_enable;
  wire  regs_383_clock;
  wire  regs_383_reset;
  wire [63:0] regs_383_io_in;
  wire [63:0] regs_383_io_init;
  wire  regs_383_io_reset;
  wire [63:0] regs_383_io_out;
  wire  regs_383_io_enable;
  wire  regs_384_clock;
  wire  regs_384_reset;
  wire [63:0] regs_384_io_in;
  wire [63:0] regs_384_io_init;
  wire  regs_384_io_reset;
  wire [63:0] regs_384_io_out;
  wire  regs_384_io_enable;
  wire  regs_385_clock;
  wire  regs_385_reset;
  wire [63:0] regs_385_io_in;
  wire [63:0] regs_385_io_init;
  wire  regs_385_io_reset;
  wire [63:0] regs_385_io_out;
  wire  regs_385_io_enable;
  wire  regs_386_clock;
  wire  regs_386_reset;
  wire [63:0] regs_386_io_in;
  wire [63:0] regs_386_io_init;
  wire  regs_386_io_reset;
  wire [63:0] regs_386_io_out;
  wire  regs_386_io_enable;
  wire  regs_387_clock;
  wire  regs_387_reset;
  wire [63:0] regs_387_io_in;
  wire [63:0] regs_387_io_init;
  wire  regs_387_io_reset;
  wire [63:0] regs_387_io_out;
  wire  regs_387_io_enable;
  wire  regs_388_clock;
  wire  regs_388_reset;
  wire [63:0] regs_388_io_in;
  wire [63:0] regs_388_io_init;
  wire  regs_388_io_reset;
  wire [63:0] regs_388_io_out;
  wire  regs_388_io_enable;
  wire  regs_389_clock;
  wire  regs_389_reset;
  wire [63:0] regs_389_io_in;
  wire [63:0] regs_389_io_init;
  wire  regs_389_io_reset;
  wire [63:0] regs_389_io_out;
  wire  regs_389_io_enable;
  wire  regs_390_clock;
  wire  regs_390_reset;
  wire [63:0] regs_390_io_in;
  wire [63:0] regs_390_io_init;
  wire  regs_390_io_reset;
  wire [63:0] regs_390_io_out;
  wire  regs_390_io_enable;
  wire  regs_391_clock;
  wire  regs_391_reset;
  wire [63:0] regs_391_io_in;
  wire [63:0] regs_391_io_init;
  wire  regs_391_io_reset;
  wire [63:0] regs_391_io_out;
  wire  regs_391_io_enable;
  wire  regs_392_clock;
  wire  regs_392_reset;
  wire [63:0] regs_392_io_in;
  wire [63:0] regs_392_io_init;
  wire  regs_392_io_reset;
  wire [63:0] regs_392_io_out;
  wire  regs_392_io_enable;
  wire  regs_393_clock;
  wire  regs_393_reset;
  wire [63:0] regs_393_io_in;
  wire [63:0] regs_393_io_init;
  wire  regs_393_io_reset;
  wire [63:0] regs_393_io_out;
  wire  regs_393_io_enable;
  wire  regs_394_clock;
  wire  regs_394_reset;
  wire [63:0] regs_394_io_in;
  wire [63:0] regs_394_io_init;
  wire  regs_394_io_reset;
  wire [63:0] regs_394_io_out;
  wire  regs_394_io_enable;
  wire  regs_395_clock;
  wire  regs_395_reset;
  wire [63:0] regs_395_io_in;
  wire [63:0] regs_395_io_init;
  wire  regs_395_io_reset;
  wire [63:0] regs_395_io_out;
  wire  regs_395_io_enable;
  wire  regs_396_clock;
  wire  regs_396_reset;
  wire [63:0] regs_396_io_in;
  wire [63:0] regs_396_io_init;
  wire  regs_396_io_reset;
  wire [63:0] regs_396_io_out;
  wire  regs_396_io_enable;
  wire  regs_397_clock;
  wire  regs_397_reset;
  wire [63:0] regs_397_io_in;
  wire [63:0] regs_397_io_init;
  wire  regs_397_io_reset;
  wire [63:0] regs_397_io_out;
  wire  regs_397_io_enable;
  wire  regs_398_clock;
  wire  regs_398_reset;
  wire [63:0] regs_398_io_in;
  wire [63:0] regs_398_io_init;
  wire  regs_398_io_reset;
  wire [63:0] regs_398_io_out;
  wire  regs_398_io_enable;
  wire  regs_399_clock;
  wire  regs_399_reset;
  wire [63:0] regs_399_io_in;
  wire [63:0] regs_399_io_init;
  wire  regs_399_io_reset;
  wire [63:0] regs_399_io_out;
  wire  regs_399_io_enable;
  wire  regs_400_clock;
  wire  regs_400_reset;
  wire [63:0] regs_400_io_in;
  wire [63:0] regs_400_io_init;
  wire  regs_400_io_reset;
  wire [63:0] regs_400_io_out;
  wire  regs_400_io_enable;
  wire  regs_401_clock;
  wire  regs_401_reset;
  wire [63:0] regs_401_io_in;
  wire [63:0] regs_401_io_init;
  wire  regs_401_io_reset;
  wire [63:0] regs_401_io_out;
  wire  regs_401_io_enable;
  wire  regs_402_clock;
  wire  regs_402_reset;
  wire [63:0] regs_402_io_in;
  wire [63:0] regs_402_io_init;
  wire  regs_402_io_reset;
  wire [63:0] regs_402_io_out;
  wire  regs_402_io_enable;
  wire  regs_403_clock;
  wire  regs_403_reset;
  wire [63:0] regs_403_io_in;
  wire [63:0] regs_403_io_init;
  wire  regs_403_io_reset;
  wire [63:0] regs_403_io_out;
  wire  regs_403_io_enable;
  wire  regs_404_clock;
  wire  regs_404_reset;
  wire [63:0] regs_404_io_in;
  wire [63:0] regs_404_io_init;
  wire  regs_404_io_reset;
  wire [63:0] regs_404_io_out;
  wire  regs_404_io_enable;
  wire  regs_405_clock;
  wire  regs_405_reset;
  wire [63:0] regs_405_io_in;
  wire [63:0] regs_405_io_init;
  wire  regs_405_io_reset;
  wire [63:0] regs_405_io_out;
  wire  regs_405_io_enable;
  wire  regs_406_clock;
  wire  regs_406_reset;
  wire [63:0] regs_406_io_in;
  wire [63:0] regs_406_io_init;
  wire  regs_406_io_reset;
  wire [63:0] regs_406_io_out;
  wire  regs_406_io_enable;
  wire  regs_407_clock;
  wire  regs_407_reset;
  wire [63:0] regs_407_io_in;
  wire [63:0] regs_407_io_init;
  wire  regs_407_io_reset;
  wire [63:0] regs_407_io_out;
  wire  regs_407_io_enable;
  wire  regs_408_clock;
  wire  regs_408_reset;
  wire [63:0] regs_408_io_in;
  wire [63:0] regs_408_io_init;
  wire  regs_408_io_reset;
  wire [63:0] regs_408_io_out;
  wire  regs_408_io_enable;
  wire  regs_409_clock;
  wire  regs_409_reset;
  wire [63:0] regs_409_io_in;
  wire [63:0] regs_409_io_init;
  wire  regs_409_io_reset;
  wire [63:0] regs_409_io_out;
  wire  regs_409_io_enable;
  wire  regs_410_clock;
  wire  regs_410_reset;
  wire [63:0] regs_410_io_in;
  wire [63:0] regs_410_io_init;
  wire  regs_410_io_reset;
  wire [63:0] regs_410_io_out;
  wire  regs_410_io_enable;
  wire  regs_411_clock;
  wire  regs_411_reset;
  wire [63:0] regs_411_io_in;
  wire [63:0] regs_411_io_init;
  wire  regs_411_io_reset;
  wire [63:0] regs_411_io_out;
  wire  regs_411_io_enable;
  wire  regs_412_clock;
  wire  regs_412_reset;
  wire [63:0] regs_412_io_in;
  wire [63:0] regs_412_io_init;
  wire  regs_412_io_reset;
  wire [63:0] regs_412_io_out;
  wire  regs_412_io_enable;
  wire  regs_413_clock;
  wire  regs_413_reset;
  wire [63:0] regs_413_io_in;
  wire [63:0] regs_413_io_init;
  wire  regs_413_io_reset;
  wire [63:0] regs_413_io_out;
  wire  regs_413_io_enable;
  wire  regs_414_clock;
  wire  regs_414_reset;
  wire [63:0] regs_414_io_in;
  wire [63:0] regs_414_io_init;
  wire  regs_414_io_reset;
  wire [63:0] regs_414_io_out;
  wire  regs_414_io_enable;
  wire  regs_415_clock;
  wire  regs_415_reset;
  wire [63:0] regs_415_io_in;
  wire [63:0] regs_415_io_init;
  wire  regs_415_io_reset;
  wire [63:0] regs_415_io_out;
  wire  regs_415_io_enable;
  wire  regs_416_clock;
  wire  regs_416_reset;
  wire [63:0] regs_416_io_in;
  wire [63:0] regs_416_io_init;
  wire  regs_416_io_reset;
  wire [63:0] regs_416_io_out;
  wire  regs_416_io_enable;
  wire  regs_417_clock;
  wire  regs_417_reset;
  wire [63:0] regs_417_io_in;
  wire [63:0] regs_417_io_init;
  wire  regs_417_io_reset;
  wire [63:0] regs_417_io_out;
  wire  regs_417_io_enable;
  wire  regs_418_clock;
  wire  regs_418_reset;
  wire [63:0] regs_418_io_in;
  wire [63:0] regs_418_io_init;
  wire  regs_418_io_reset;
  wire [63:0] regs_418_io_out;
  wire  regs_418_io_enable;
  wire  regs_419_clock;
  wire  regs_419_reset;
  wire [63:0] regs_419_io_in;
  wire [63:0] regs_419_io_init;
  wire  regs_419_io_reset;
  wire [63:0] regs_419_io_out;
  wire  regs_419_io_enable;
  wire  regs_420_clock;
  wire  regs_420_reset;
  wire [63:0] regs_420_io_in;
  wire [63:0] regs_420_io_init;
  wire  regs_420_io_reset;
  wire [63:0] regs_420_io_out;
  wire  regs_420_io_enable;
  wire  regs_421_clock;
  wire  regs_421_reset;
  wire [63:0] regs_421_io_in;
  wire [63:0] regs_421_io_init;
  wire  regs_421_io_reset;
  wire [63:0] regs_421_io_out;
  wire  regs_421_io_enable;
  wire  regs_422_clock;
  wire  regs_422_reset;
  wire [63:0] regs_422_io_in;
  wire [63:0] regs_422_io_init;
  wire  regs_422_io_reset;
  wire [63:0] regs_422_io_out;
  wire  regs_422_io_enable;
  wire  regs_423_clock;
  wire  regs_423_reset;
  wire [63:0] regs_423_io_in;
  wire [63:0] regs_423_io_init;
  wire  regs_423_io_reset;
  wire [63:0] regs_423_io_out;
  wire  regs_423_io_enable;
  wire  regs_424_clock;
  wire  regs_424_reset;
  wire [63:0] regs_424_io_in;
  wire [63:0] regs_424_io_init;
  wire  regs_424_io_reset;
  wire [63:0] regs_424_io_out;
  wire  regs_424_io_enable;
  wire  regs_425_clock;
  wire  regs_425_reset;
  wire [63:0] regs_425_io_in;
  wire [63:0] regs_425_io_init;
  wire  regs_425_io_reset;
  wire [63:0] regs_425_io_out;
  wire  regs_425_io_enable;
  wire  regs_426_clock;
  wire  regs_426_reset;
  wire [63:0] regs_426_io_in;
  wire [63:0] regs_426_io_init;
  wire  regs_426_io_reset;
  wire [63:0] regs_426_io_out;
  wire  regs_426_io_enable;
  wire  regs_427_clock;
  wire  regs_427_reset;
  wire [63:0] regs_427_io_in;
  wire [63:0] regs_427_io_init;
  wire  regs_427_io_reset;
  wire [63:0] regs_427_io_out;
  wire  regs_427_io_enable;
  wire  regs_428_clock;
  wire  regs_428_reset;
  wire [63:0] regs_428_io_in;
  wire [63:0] regs_428_io_init;
  wire  regs_428_io_reset;
  wire [63:0] regs_428_io_out;
  wire  regs_428_io_enable;
  wire  regs_429_clock;
  wire  regs_429_reset;
  wire [63:0] regs_429_io_in;
  wire [63:0] regs_429_io_init;
  wire  regs_429_io_reset;
  wire [63:0] regs_429_io_out;
  wire  regs_429_io_enable;
  wire  regs_430_clock;
  wire  regs_430_reset;
  wire [63:0] regs_430_io_in;
  wire [63:0] regs_430_io_init;
  wire  regs_430_io_reset;
  wire [63:0] regs_430_io_out;
  wire  regs_430_io_enable;
  wire  regs_431_clock;
  wire  regs_431_reset;
  wire [63:0] regs_431_io_in;
  wire [63:0] regs_431_io_init;
  wire  regs_431_io_reset;
  wire [63:0] regs_431_io_out;
  wire  regs_431_io_enable;
  wire  regs_432_clock;
  wire  regs_432_reset;
  wire [63:0] regs_432_io_in;
  wire [63:0] regs_432_io_init;
  wire  regs_432_io_reset;
  wire [63:0] regs_432_io_out;
  wire  regs_432_io_enable;
  wire  regs_433_clock;
  wire  regs_433_reset;
  wire [63:0] regs_433_io_in;
  wire [63:0] regs_433_io_init;
  wire  regs_433_io_reset;
  wire [63:0] regs_433_io_out;
  wire  regs_433_io_enable;
  wire  regs_434_clock;
  wire  regs_434_reset;
  wire [63:0] regs_434_io_in;
  wire [63:0] regs_434_io_init;
  wire  regs_434_io_reset;
  wire [63:0] regs_434_io_out;
  wire  regs_434_io_enable;
  wire  regs_435_clock;
  wire  regs_435_reset;
  wire [63:0] regs_435_io_in;
  wire [63:0] regs_435_io_init;
  wire  regs_435_io_reset;
  wire [63:0] regs_435_io_out;
  wire  regs_435_io_enable;
  wire  regs_436_clock;
  wire  regs_436_reset;
  wire [63:0] regs_436_io_in;
  wire [63:0] regs_436_io_init;
  wire  regs_436_io_reset;
  wire [63:0] regs_436_io_out;
  wire  regs_436_io_enable;
  wire  regs_437_clock;
  wire  regs_437_reset;
  wire [63:0] regs_437_io_in;
  wire [63:0] regs_437_io_init;
  wire  regs_437_io_reset;
  wire [63:0] regs_437_io_out;
  wire  regs_437_io_enable;
  wire  regs_438_clock;
  wire  regs_438_reset;
  wire [63:0] regs_438_io_in;
  wire [63:0] regs_438_io_init;
  wire  regs_438_io_reset;
  wire [63:0] regs_438_io_out;
  wire  regs_438_io_enable;
  wire  regs_439_clock;
  wire  regs_439_reset;
  wire [63:0] regs_439_io_in;
  wire [63:0] regs_439_io_init;
  wire  regs_439_io_reset;
  wire [63:0] regs_439_io_out;
  wire  regs_439_io_enable;
  wire  regs_440_clock;
  wire  regs_440_reset;
  wire [63:0] regs_440_io_in;
  wire [63:0] regs_440_io_init;
  wire  regs_440_io_reset;
  wire [63:0] regs_440_io_out;
  wire  regs_440_io_enable;
  wire  regs_441_clock;
  wire  regs_441_reset;
  wire [63:0] regs_441_io_in;
  wire [63:0] regs_441_io_init;
  wire  regs_441_io_reset;
  wire [63:0] regs_441_io_out;
  wire  regs_441_io_enable;
  wire  regs_442_clock;
  wire  regs_442_reset;
  wire [63:0] regs_442_io_in;
  wire [63:0] regs_442_io_init;
  wire  regs_442_io_reset;
  wire [63:0] regs_442_io_out;
  wire  regs_442_io_enable;
  wire  regs_443_clock;
  wire  regs_443_reset;
  wire [63:0] regs_443_io_in;
  wire [63:0] regs_443_io_init;
  wire  regs_443_io_reset;
  wire [63:0] regs_443_io_out;
  wire  regs_443_io_enable;
  wire  regs_444_clock;
  wire  regs_444_reset;
  wire [63:0] regs_444_io_in;
  wire [63:0] regs_444_io_init;
  wire  regs_444_io_reset;
  wire [63:0] regs_444_io_out;
  wire  regs_444_io_enable;
  wire  regs_445_clock;
  wire  regs_445_reset;
  wire [63:0] regs_445_io_in;
  wire [63:0] regs_445_io_init;
  wire  regs_445_io_reset;
  wire [63:0] regs_445_io_out;
  wire  regs_445_io_enable;
  wire  regs_446_clock;
  wire  regs_446_reset;
  wire [63:0] regs_446_io_in;
  wire [63:0] regs_446_io_init;
  wire  regs_446_io_reset;
  wire [63:0] regs_446_io_out;
  wire  regs_446_io_enable;
  wire  regs_447_clock;
  wire  regs_447_reset;
  wire [63:0] regs_447_io_in;
  wire [63:0] regs_447_io_init;
  wire  regs_447_io_reset;
  wire [63:0] regs_447_io_out;
  wire  regs_447_io_enable;
  wire  regs_448_clock;
  wire  regs_448_reset;
  wire [63:0] regs_448_io_in;
  wire [63:0] regs_448_io_init;
  wire  regs_448_io_reset;
  wire [63:0] regs_448_io_out;
  wire  regs_448_io_enable;
  wire  regs_449_clock;
  wire  regs_449_reset;
  wire [63:0] regs_449_io_in;
  wire [63:0] regs_449_io_init;
  wire  regs_449_io_reset;
  wire [63:0] regs_449_io_out;
  wire  regs_449_io_enable;
  wire  regs_450_clock;
  wire  regs_450_reset;
  wire [63:0] regs_450_io_in;
  wire [63:0] regs_450_io_init;
  wire  regs_450_io_reset;
  wire [63:0] regs_450_io_out;
  wire  regs_450_io_enable;
  wire  regs_451_clock;
  wire  regs_451_reset;
  wire [63:0] regs_451_io_in;
  wire [63:0] regs_451_io_init;
  wire  regs_451_io_reset;
  wire [63:0] regs_451_io_out;
  wire  regs_451_io_enable;
  wire  regs_452_clock;
  wire  regs_452_reset;
  wire [63:0] regs_452_io_in;
  wire [63:0] regs_452_io_init;
  wire  regs_452_io_reset;
  wire [63:0] regs_452_io_out;
  wire  regs_452_io_enable;
  wire  regs_453_clock;
  wire  regs_453_reset;
  wire [63:0] regs_453_io_in;
  wire [63:0] regs_453_io_init;
  wire  regs_453_io_reset;
  wire [63:0] regs_453_io_out;
  wire  regs_453_io_enable;
  wire  regs_454_clock;
  wire  regs_454_reset;
  wire [63:0] regs_454_io_in;
  wire [63:0] regs_454_io_init;
  wire  regs_454_io_reset;
  wire [63:0] regs_454_io_out;
  wire  regs_454_io_enable;
  wire  regs_455_clock;
  wire  regs_455_reset;
  wire [63:0] regs_455_io_in;
  wire [63:0] regs_455_io_init;
  wire  regs_455_io_reset;
  wire [63:0] regs_455_io_out;
  wire  regs_455_io_enable;
  wire  regs_456_clock;
  wire  regs_456_reset;
  wire [63:0] regs_456_io_in;
  wire [63:0] regs_456_io_init;
  wire  regs_456_io_reset;
  wire [63:0] regs_456_io_out;
  wire  regs_456_io_enable;
  wire  regs_457_clock;
  wire  regs_457_reset;
  wire [63:0] regs_457_io_in;
  wire [63:0] regs_457_io_init;
  wire  regs_457_io_reset;
  wire [63:0] regs_457_io_out;
  wire  regs_457_io_enable;
  wire  regs_458_clock;
  wire  regs_458_reset;
  wire [63:0] regs_458_io_in;
  wire [63:0] regs_458_io_init;
  wire  regs_458_io_reset;
  wire [63:0] regs_458_io_out;
  wire  regs_458_io_enable;
  wire  regs_459_clock;
  wire  regs_459_reset;
  wire [63:0] regs_459_io_in;
  wire [63:0] regs_459_io_init;
  wire  regs_459_io_reset;
  wire [63:0] regs_459_io_out;
  wire  regs_459_io_enable;
  wire  regs_460_clock;
  wire  regs_460_reset;
  wire [63:0] regs_460_io_in;
  wire [63:0] regs_460_io_init;
  wire  regs_460_io_reset;
  wire [63:0] regs_460_io_out;
  wire  regs_460_io_enable;
  wire  regs_461_clock;
  wire  regs_461_reset;
  wire [63:0] regs_461_io_in;
  wire [63:0] regs_461_io_init;
  wire  regs_461_io_reset;
  wire [63:0] regs_461_io_out;
  wire  regs_461_io_enable;
  wire  regs_462_clock;
  wire  regs_462_reset;
  wire [63:0] regs_462_io_in;
  wire [63:0] regs_462_io_init;
  wire  regs_462_io_reset;
  wire [63:0] regs_462_io_out;
  wire  regs_462_io_enable;
  wire  regs_463_clock;
  wire  regs_463_reset;
  wire [63:0] regs_463_io_in;
  wire [63:0] regs_463_io_init;
  wire  regs_463_io_reset;
  wire [63:0] regs_463_io_out;
  wire  regs_463_io_enable;
  wire  regs_464_clock;
  wire  regs_464_reset;
  wire [63:0] regs_464_io_in;
  wire [63:0] regs_464_io_init;
  wire  regs_464_io_reset;
  wire [63:0] regs_464_io_out;
  wire  regs_464_io_enable;
  wire  regs_465_clock;
  wire  regs_465_reset;
  wire [63:0] regs_465_io_in;
  wire [63:0] regs_465_io_init;
  wire  regs_465_io_reset;
  wire [63:0] regs_465_io_out;
  wire  regs_465_io_enable;
  wire  regs_466_clock;
  wire  regs_466_reset;
  wire [63:0] regs_466_io_in;
  wire [63:0] regs_466_io_init;
  wire  regs_466_io_reset;
  wire [63:0] regs_466_io_out;
  wire  regs_466_io_enable;
  wire  regs_467_clock;
  wire  regs_467_reset;
  wire [63:0] regs_467_io_in;
  wire [63:0] regs_467_io_init;
  wire  regs_467_io_reset;
  wire [63:0] regs_467_io_out;
  wire  regs_467_io_enable;
  wire  regs_468_clock;
  wire  regs_468_reset;
  wire [63:0] regs_468_io_in;
  wire [63:0] regs_468_io_init;
  wire  regs_468_io_reset;
  wire [63:0] regs_468_io_out;
  wire  regs_468_io_enable;
  wire  regs_469_clock;
  wire  regs_469_reset;
  wire [63:0] regs_469_io_in;
  wire [63:0] regs_469_io_init;
  wire  regs_469_io_reset;
  wire [63:0] regs_469_io_out;
  wire  regs_469_io_enable;
  wire  regs_470_clock;
  wire  regs_470_reset;
  wire [63:0] regs_470_io_in;
  wire [63:0] regs_470_io_init;
  wire  regs_470_io_reset;
  wire [63:0] regs_470_io_out;
  wire  regs_470_io_enable;
  wire  regs_471_clock;
  wire  regs_471_reset;
  wire [63:0] regs_471_io_in;
  wire [63:0] regs_471_io_init;
  wire  regs_471_io_reset;
  wire [63:0] regs_471_io_out;
  wire  regs_471_io_enable;
  wire  regs_472_clock;
  wire  regs_472_reset;
  wire [63:0] regs_472_io_in;
  wire [63:0] regs_472_io_init;
  wire  regs_472_io_reset;
  wire [63:0] regs_472_io_out;
  wire  regs_472_io_enable;
  wire  regs_473_clock;
  wire  regs_473_reset;
  wire [63:0] regs_473_io_in;
  wire [63:0] regs_473_io_init;
  wire  regs_473_io_reset;
  wire [63:0] regs_473_io_out;
  wire  regs_473_io_enable;
  wire  regs_474_clock;
  wire  regs_474_reset;
  wire [63:0] regs_474_io_in;
  wire [63:0] regs_474_io_init;
  wire  regs_474_io_reset;
  wire [63:0] regs_474_io_out;
  wire  regs_474_io_enable;
  wire  regs_475_clock;
  wire  regs_475_reset;
  wire [63:0] regs_475_io_in;
  wire [63:0] regs_475_io_init;
  wire  regs_475_io_reset;
  wire [63:0] regs_475_io_out;
  wire  regs_475_io_enable;
  wire  regs_476_clock;
  wire  regs_476_reset;
  wire [63:0] regs_476_io_in;
  wire [63:0] regs_476_io_init;
  wire  regs_476_io_reset;
  wire [63:0] regs_476_io_out;
  wire  regs_476_io_enable;
  wire  regs_477_clock;
  wire  regs_477_reset;
  wire [63:0] regs_477_io_in;
  wire [63:0] regs_477_io_init;
  wire  regs_477_io_reset;
  wire [63:0] regs_477_io_out;
  wire  regs_477_io_enable;
  wire  regs_478_clock;
  wire  regs_478_reset;
  wire [63:0] regs_478_io_in;
  wire [63:0] regs_478_io_init;
  wire  regs_478_io_reset;
  wire [63:0] regs_478_io_out;
  wire  regs_478_io_enable;
  wire  regs_479_clock;
  wire  regs_479_reset;
  wire [63:0] regs_479_io_in;
  wire [63:0] regs_479_io_init;
  wire  regs_479_io_reset;
  wire [63:0] regs_479_io_out;
  wire  regs_479_io_enable;
  wire  regs_480_clock;
  wire  regs_480_reset;
  wire [63:0] regs_480_io_in;
  wire [63:0] regs_480_io_init;
  wire  regs_480_io_reset;
  wire [63:0] regs_480_io_out;
  wire  regs_480_io_enable;
  wire  regs_481_clock;
  wire  regs_481_reset;
  wire [63:0] regs_481_io_in;
  wire [63:0] regs_481_io_init;
  wire  regs_481_io_reset;
  wire [63:0] regs_481_io_out;
  wire  regs_481_io_enable;
  wire  regs_482_clock;
  wire  regs_482_reset;
  wire [63:0] regs_482_io_in;
  wire [63:0] regs_482_io_init;
  wire  regs_482_io_reset;
  wire [63:0] regs_482_io_out;
  wire  regs_482_io_enable;
  wire  regs_483_clock;
  wire  regs_483_reset;
  wire [63:0] regs_483_io_in;
  wire [63:0] regs_483_io_init;
  wire  regs_483_io_reset;
  wire [63:0] regs_483_io_out;
  wire  regs_483_io_enable;
  wire  regs_484_clock;
  wire  regs_484_reset;
  wire [63:0] regs_484_io_in;
  wire [63:0] regs_484_io_init;
  wire  regs_484_io_reset;
  wire [63:0] regs_484_io_out;
  wire  regs_484_io_enable;
  wire  regs_485_clock;
  wire  regs_485_reset;
  wire [63:0] regs_485_io_in;
  wire [63:0] regs_485_io_init;
  wire  regs_485_io_reset;
  wire [63:0] regs_485_io_out;
  wire  regs_485_io_enable;
  wire  regs_486_clock;
  wire  regs_486_reset;
  wire [63:0] regs_486_io_in;
  wire [63:0] regs_486_io_init;
  wire  regs_486_io_reset;
  wire [63:0] regs_486_io_out;
  wire  regs_486_io_enable;
  wire  regs_487_clock;
  wire  regs_487_reset;
  wire [63:0] regs_487_io_in;
  wire [63:0] regs_487_io_init;
  wire  regs_487_io_reset;
  wire [63:0] regs_487_io_out;
  wire  regs_487_io_enable;
  wire  regs_488_clock;
  wire  regs_488_reset;
  wire [63:0] regs_488_io_in;
  wire [63:0] regs_488_io_init;
  wire  regs_488_io_reset;
  wire [63:0] regs_488_io_out;
  wire  regs_488_io_enable;
  wire  regs_489_clock;
  wire  regs_489_reset;
  wire [63:0] regs_489_io_in;
  wire [63:0] regs_489_io_init;
  wire  regs_489_io_reset;
  wire [63:0] regs_489_io_out;
  wire  regs_489_io_enable;
  wire  regs_490_clock;
  wire  regs_490_reset;
  wire [63:0] regs_490_io_in;
  wire [63:0] regs_490_io_init;
  wire  regs_490_io_reset;
  wire [63:0] regs_490_io_out;
  wire  regs_490_io_enable;
  wire  regs_491_clock;
  wire  regs_491_reset;
  wire [63:0] regs_491_io_in;
  wire [63:0] regs_491_io_init;
  wire  regs_491_io_reset;
  wire [63:0] regs_491_io_out;
  wire  regs_491_io_enable;
  wire  regs_492_clock;
  wire  regs_492_reset;
  wire [63:0] regs_492_io_in;
  wire [63:0] regs_492_io_init;
  wire  regs_492_io_reset;
  wire [63:0] regs_492_io_out;
  wire  regs_492_io_enable;
  wire  regs_493_clock;
  wire  regs_493_reset;
  wire [63:0] regs_493_io_in;
  wire [63:0] regs_493_io_init;
  wire  regs_493_io_reset;
  wire [63:0] regs_493_io_out;
  wire  regs_493_io_enable;
  wire  regs_494_clock;
  wire  regs_494_reset;
  wire [63:0] regs_494_io_in;
  wire [63:0] regs_494_io_init;
  wire  regs_494_io_reset;
  wire [63:0] regs_494_io_out;
  wire  regs_494_io_enable;
  wire  regs_495_clock;
  wire  regs_495_reset;
  wire [63:0] regs_495_io_in;
  wire [63:0] regs_495_io_init;
  wire  regs_495_io_reset;
  wire [63:0] regs_495_io_out;
  wire  regs_495_io_enable;
  wire  regs_496_clock;
  wire  regs_496_reset;
  wire [63:0] regs_496_io_in;
  wire [63:0] regs_496_io_init;
  wire  regs_496_io_reset;
  wire [63:0] regs_496_io_out;
  wire  regs_496_io_enable;
  wire  regs_497_clock;
  wire  regs_497_reset;
  wire [63:0] regs_497_io_in;
  wire [63:0] regs_497_io_init;
  wire  regs_497_io_reset;
  wire [63:0] regs_497_io_out;
  wire  regs_497_io_enable;
  wire  regs_498_clock;
  wire  regs_498_reset;
  wire [63:0] regs_498_io_in;
  wire [63:0] regs_498_io_init;
  wire  regs_498_io_reset;
  wire [63:0] regs_498_io_out;
  wire  regs_498_io_enable;
  wire  regs_499_clock;
  wire  regs_499_reset;
  wire [63:0] regs_499_io_in;
  wire [63:0] regs_499_io_init;
  wire  regs_499_io_reset;
  wire [63:0] regs_499_io_out;
  wire  regs_499_io_enable;
  wire  regs_500_clock;
  wire  regs_500_reset;
  wire [63:0] regs_500_io_in;
  wire [63:0] regs_500_io_init;
  wire  regs_500_io_reset;
  wire [63:0] regs_500_io_out;
  wire  regs_500_io_enable;
  wire  regs_501_clock;
  wire  regs_501_reset;
  wire [63:0] regs_501_io_in;
  wire [63:0] regs_501_io_init;
  wire  regs_501_io_reset;
  wire [63:0] regs_501_io_out;
  wire  regs_501_io_enable;
  wire  regs_502_clock;
  wire  regs_502_reset;
  wire [63:0] regs_502_io_in;
  wire [63:0] regs_502_io_init;
  wire  regs_502_io_reset;
  wire [63:0] regs_502_io_out;
  wire  regs_502_io_enable;
  wire  regs_503_clock;
  wire  regs_503_reset;
  wire [63:0] regs_503_io_in;
  wire [63:0] regs_503_io_init;
  wire  regs_503_io_reset;
  wire [63:0] regs_503_io_out;
  wire  regs_503_io_enable;
  wire  regs_504_clock;
  wire  regs_504_reset;
  wire [63:0] regs_504_io_in;
  wire [63:0] regs_504_io_init;
  wire  regs_504_io_reset;
  wire [63:0] regs_504_io_out;
  wire  regs_504_io_enable;
  wire  regs_505_clock;
  wire  regs_505_reset;
  wire [63:0] regs_505_io_in;
  wire [63:0] regs_505_io_init;
  wire  regs_505_io_reset;
  wire [63:0] regs_505_io_out;
  wire  regs_505_io_enable;
  wire [63:0] rport_io_ins_0;
  wire [63:0] rport_io_ins_1;
  wire [63:0] rport_io_ins_2;
  wire [63:0] rport_io_ins_3;
  wire [63:0] rport_io_ins_4;
  wire [63:0] rport_io_ins_5;
  wire [63:0] rport_io_ins_6;
  wire [63:0] rport_io_ins_7;
  wire [63:0] rport_io_ins_8;
  wire [63:0] rport_io_ins_9;
  wire [63:0] rport_io_ins_10;
  wire [63:0] rport_io_ins_11;
  wire [63:0] rport_io_ins_12;
  wire [63:0] rport_io_ins_13;
  wire [63:0] rport_io_ins_14;
  wire [63:0] rport_io_ins_15;
  wire [63:0] rport_io_ins_16;
  wire [63:0] rport_io_ins_17;
  wire [63:0] rport_io_ins_18;
  wire [63:0] rport_io_ins_19;
  wire [63:0] rport_io_ins_20;
  wire [63:0] rport_io_ins_21;
  wire [63:0] rport_io_ins_22;
  wire [63:0] rport_io_ins_23;
  wire [63:0] rport_io_ins_24;
  wire [63:0] rport_io_ins_25;
  wire [63:0] rport_io_ins_26;
  wire [63:0] rport_io_ins_27;
  wire [63:0] rport_io_ins_28;
  wire [63:0] rport_io_ins_29;
  wire [63:0] rport_io_ins_30;
  wire [63:0] rport_io_ins_31;
  wire [63:0] rport_io_ins_32;
  wire [63:0] rport_io_ins_33;
  wire [63:0] rport_io_ins_34;
  wire [63:0] rport_io_ins_35;
  wire [63:0] rport_io_ins_36;
  wire [63:0] rport_io_ins_37;
  wire [63:0] rport_io_ins_38;
  wire [63:0] rport_io_ins_39;
  wire [63:0] rport_io_ins_40;
  wire [63:0] rport_io_ins_41;
  wire [63:0] rport_io_ins_42;
  wire [63:0] rport_io_ins_43;
  wire [63:0] rport_io_ins_44;
  wire [63:0] rport_io_ins_45;
  wire [63:0] rport_io_ins_46;
  wire [63:0] rport_io_ins_47;
  wire [63:0] rport_io_ins_48;
  wire [63:0] rport_io_ins_49;
  wire [63:0] rport_io_ins_50;
  wire [63:0] rport_io_ins_51;
  wire [63:0] rport_io_ins_52;
  wire [63:0] rport_io_ins_53;
  wire [63:0] rport_io_ins_54;
  wire [63:0] rport_io_ins_55;
  wire [63:0] rport_io_ins_56;
  wire [63:0] rport_io_ins_57;
  wire [63:0] rport_io_ins_58;
  wire [63:0] rport_io_ins_59;
  wire [63:0] rport_io_ins_60;
  wire [63:0] rport_io_ins_61;
  wire [63:0] rport_io_ins_62;
  wire [63:0] rport_io_ins_63;
  wire [63:0] rport_io_ins_64;
  wire [63:0] rport_io_ins_65;
  wire [63:0] rport_io_ins_66;
  wire [63:0] rport_io_ins_67;
  wire [63:0] rport_io_ins_68;
  wire [63:0] rport_io_ins_69;
  wire [63:0] rport_io_ins_70;
  wire [63:0] rport_io_ins_71;
  wire [63:0] rport_io_ins_72;
  wire [63:0] rport_io_ins_73;
  wire [63:0] rport_io_ins_74;
  wire [63:0] rport_io_ins_75;
  wire [63:0] rport_io_ins_76;
  wire [63:0] rport_io_ins_77;
  wire [63:0] rport_io_ins_78;
  wire [63:0] rport_io_ins_79;
  wire [63:0] rport_io_ins_80;
  wire [63:0] rport_io_ins_81;
  wire [63:0] rport_io_ins_82;
  wire [63:0] rport_io_ins_83;
  wire [63:0] rport_io_ins_84;
  wire [63:0] rport_io_ins_85;
  wire [63:0] rport_io_ins_86;
  wire [63:0] rport_io_ins_87;
  wire [63:0] rport_io_ins_88;
  wire [63:0] rport_io_ins_89;
  wire [63:0] rport_io_ins_90;
  wire [63:0] rport_io_ins_91;
  wire [63:0] rport_io_ins_92;
  wire [63:0] rport_io_ins_93;
  wire [63:0] rport_io_ins_94;
  wire [63:0] rport_io_ins_95;
  wire [63:0] rport_io_ins_96;
  wire [63:0] rport_io_ins_97;
  wire [63:0] rport_io_ins_98;
  wire [63:0] rport_io_ins_99;
  wire [63:0] rport_io_ins_100;
  wire [63:0] rport_io_ins_101;
  wire [63:0] rport_io_ins_102;
  wire [63:0] rport_io_ins_103;
  wire [63:0] rport_io_ins_104;
  wire [63:0] rport_io_ins_105;
  wire [63:0] rport_io_ins_106;
  wire [63:0] rport_io_ins_107;
  wire [63:0] rport_io_ins_108;
  wire [63:0] rport_io_ins_109;
  wire [63:0] rport_io_ins_110;
  wire [63:0] rport_io_ins_111;
  wire [63:0] rport_io_ins_112;
  wire [63:0] rport_io_ins_113;
  wire [63:0] rport_io_ins_114;
  wire [63:0] rport_io_ins_115;
  wire [63:0] rport_io_ins_116;
  wire [63:0] rport_io_ins_117;
  wire [63:0] rport_io_ins_118;
  wire [63:0] rport_io_ins_119;
  wire [63:0] rport_io_ins_120;
  wire [63:0] rport_io_ins_121;
  wire [63:0] rport_io_ins_122;
  wire [63:0] rport_io_ins_123;
  wire [63:0] rport_io_ins_124;
  wire [63:0] rport_io_ins_125;
  wire [63:0] rport_io_ins_126;
  wire [63:0] rport_io_ins_127;
  wire [63:0] rport_io_ins_128;
  wire [63:0] rport_io_ins_129;
  wire [63:0] rport_io_ins_130;
  wire [63:0] rport_io_ins_131;
  wire [63:0] rport_io_ins_132;
  wire [63:0] rport_io_ins_133;
  wire [63:0] rport_io_ins_134;
  wire [63:0] rport_io_ins_135;
  wire [63:0] rport_io_ins_136;
  wire [63:0] rport_io_ins_137;
  wire [63:0] rport_io_ins_138;
  wire [63:0] rport_io_ins_139;
  wire [63:0] rport_io_ins_140;
  wire [63:0] rport_io_ins_141;
  wire [63:0] rport_io_ins_142;
  wire [63:0] rport_io_ins_143;
  wire [63:0] rport_io_ins_144;
  wire [63:0] rport_io_ins_145;
  wire [63:0] rport_io_ins_146;
  wire [63:0] rport_io_ins_147;
  wire [63:0] rport_io_ins_148;
  wire [63:0] rport_io_ins_149;
  wire [63:0] rport_io_ins_150;
  wire [63:0] rport_io_ins_151;
  wire [63:0] rport_io_ins_152;
  wire [63:0] rport_io_ins_153;
  wire [63:0] rport_io_ins_154;
  wire [63:0] rport_io_ins_155;
  wire [63:0] rport_io_ins_156;
  wire [63:0] rport_io_ins_157;
  wire [63:0] rport_io_ins_158;
  wire [63:0] rport_io_ins_159;
  wire [63:0] rport_io_ins_160;
  wire [63:0] rport_io_ins_161;
  wire [63:0] rport_io_ins_162;
  wire [63:0] rport_io_ins_163;
  wire [63:0] rport_io_ins_164;
  wire [63:0] rport_io_ins_165;
  wire [63:0] rport_io_ins_166;
  wire [63:0] rport_io_ins_167;
  wire [63:0] rport_io_ins_168;
  wire [63:0] rport_io_ins_169;
  wire [63:0] rport_io_ins_170;
  wire [63:0] rport_io_ins_171;
  wire [63:0] rport_io_ins_172;
  wire [63:0] rport_io_ins_173;
  wire [63:0] rport_io_ins_174;
  wire [63:0] rport_io_ins_175;
  wire [63:0] rport_io_ins_176;
  wire [63:0] rport_io_ins_177;
  wire [63:0] rport_io_ins_178;
  wire [63:0] rport_io_ins_179;
  wire [63:0] rport_io_ins_180;
  wire [63:0] rport_io_ins_181;
  wire [63:0] rport_io_ins_182;
  wire [63:0] rport_io_ins_183;
  wire [63:0] rport_io_ins_184;
  wire [63:0] rport_io_ins_185;
  wire [63:0] rport_io_ins_186;
  wire [63:0] rport_io_ins_187;
  wire [63:0] rport_io_ins_188;
  wire [63:0] rport_io_ins_189;
  wire [63:0] rport_io_ins_190;
  wire [63:0] rport_io_ins_191;
  wire [63:0] rport_io_ins_192;
  wire [63:0] rport_io_ins_193;
  wire [63:0] rport_io_ins_194;
  wire [63:0] rport_io_ins_195;
  wire [63:0] rport_io_ins_196;
  wire [63:0] rport_io_ins_197;
  wire [63:0] rport_io_ins_198;
  wire [63:0] rport_io_ins_199;
  wire [63:0] rport_io_ins_200;
  wire [63:0] rport_io_ins_201;
  wire [63:0] rport_io_ins_202;
  wire [63:0] rport_io_ins_203;
  wire [63:0] rport_io_ins_204;
  wire [63:0] rport_io_ins_205;
  wire [63:0] rport_io_ins_206;
  wire [63:0] rport_io_ins_207;
  wire [63:0] rport_io_ins_208;
  wire [63:0] rport_io_ins_209;
  wire [63:0] rport_io_ins_210;
  wire [63:0] rport_io_ins_211;
  wire [63:0] rport_io_ins_212;
  wire [63:0] rport_io_ins_213;
  wire [63:0] rport_io_ins_214;
  wire [63:0] rport_io_ins_215;
  wire [63:0] rport_io_ins_216;
  wire [63:0] rport_io_ins_217;
  wire [63:0] rport_io_ins_218;
  wire [63:0] rport_io_ins_219;
  wire [63:0] rport_io_ins_220;
  wire [63:0] rport_io_ins_221;
  wire [63:0] rport_io_ins_222;
  wire [63:0] rport_io_ins_223;
  wire [63:0] rport_io_ins_224;
  wire [63:0] rport_io_ins_225;
  wire [63:0] rport_io_ins_226;
  wire [63:0] rport_io_ins_227;
  wire [63:0] rport_io_ins_228;
  wire [63:0] rport_io_ins_229;
  wire [63:0] rport_io_ins_230;
  wire [63:0] rport_io_ins_231;
  wire [63:0] rport_io_ins_232;
  wire [63:0] rport_io_ins_233;
  wire [63:0] rport_io_ins_234;
  wire [63:0] rport_io_ins_235;
  wire [63:0] rport_io_ins_236;
  wire [63:0] rport_io_ins_237;
  wire [63:0] rport_io_ins_238;
  wire [63:0] rport_io_ins_239;
  wire [63:0] rport_io_ins_240;
  wire [63:0] rport_io_ins_241;
  wire [63:0] rport_io_ins_242;
  wire [63:0] rport_io_ins_243;
  wire [63:0] rport_io_ins_244;
  wire [63:0] rport_io_ins_245;
  wire [63:0] rport_io_ins_246;
  wire [63:0] rport_io_ins_247;
  wire [63:0] rport_io_ins_248;
  wire [63:0] rport_io_ins_249;
  wire [63:0] rport_io_ins_250;
  wire [63:0] rport_io_ins_251;
  wire [63:0] rport_io_ins_252;
  wire [63:0] rport_io_ins_253;
  wire [63:0] rport_io_ins_254;
  wire [63:0] rport_io_ins_255;
  wire [63:0] rport_io_ins_256;
  wire [63:0] rport_io_ins_257;
  wire [63:0] rport_io_ins_258;
  wire [63:0] rport_io_ins_259;
  wire [63:0] rport_io_ins_260;
  wire [63:0] rport_io_ins_261;
  wire [63:0] rport_io_ins_262;
  wire [63:0] rport_io_ins_263;
  wire [63:0] rport_io_ins_264;
  wire [63:0] rport_io_ins_265;
  wire [63:0] rport_io_ins_266;
  wire [63:0] rport_io_ins_267;
  wire [63:0] rport_io_ins_268;
  wire [63:0] rport_io_ins_269;
  wire [63:0] rport_io_ins_270;
  wire [63:0] rport_io_ins_271;
  wire [63:0] rport_io_ins_272;
  wire [63:0] rport_io_ins_273;
  wire [63:0] rport_io_ins_274;
  wire [63:0] rport_io_ins_275;
  wire [63:0] rport_io_ins_276;
  wire [63:0] rport_io_ins_277;
  wire [63:0] rport_io_ins_278;
  wire [63:0] rport_io_ins_279;
  wire [63:0] rport_io_ins_280;
  wire [63:0] rport_io_ins_281;
  wire [63:0] rport_io_ins_282;
  wire [63:0] rport_io_ins_283;
  wire [63:0] rport_io_ins_284;
  wire [63:0] rport_io_ins_285;
  wire [63:0] rport_io_ins_286;
  wire [63:0] rport_io_ins_287;
  wire [63:0] rport_io_ins_288;
  wire [63:0] rport_io_ins_289;
  wire [63:0] rport_io_ins_290;
  wire [63:0] rport_io_ins_291;
  wire [63:0] rport_io_ins_292;
  wire [63:0] rport_io_ins_293;
  wire [63:0] rport_io_ins_294;
  wire [63:0] rport_io_ins_295;
  wire [63:0] rport_io_ins_296;
  wire [63:0] rport_io_ins_297;
  wire [63:0] rport_io_ins_298;
  wire [63:0] rport_io_ins_299;
  wire [63:0] rport_io_ins_300;
  wire [63:0] rport_io_ins_301;
  wire [63:0] rport_io_ins_302;
  wire [63:0] rport_io_ins_303;
  wire [63:0] rport_io_ins_304;
  wire [63:0] rport_io_ins_305;
  wire [63:0] rport_io_ins_306;
  wire [63:0] rport_io_ins_307;
  wire [63:0] rport_io_ins_308;
  wire [63:0] rport_io_ins_309;
  wire [63:0] rport_io_ins_310;
  wire [63:0] rport_io_ins_311;
  wire [63:0] rport_io_ins_312;
  wire [63:0] rport_io_ins_313;
  wire [63:0] rport_io_ins_314;
  wire [63:0] rport_io_ins_315;
  wire [63:0] rport_io_ins_316;
  wire [63:0] rport_io_ins_317;
  wire [63:0] rport_io_ins_318;
  wire [63:0] rport_io_ins_319;
  wire [63:0] rport_io_ins_320;
  wire [63:0] rport_io_ins_321;
  wire [63:0] rport_io_ins_322;
  wire [63:0] rport_io_ins_323;
  wire [63:0] rport_io_ins_324;
  wire [63:0] rport_io_ins_325;
  wire [63:0] rport_io_ins_326;
  wire [63:0] rport_io_ins_327;
  wire [63:0] rport_io_ins_328;
  wire [63:0] rport_io_ins_329;
  wire [63:0] rport_io_ins_330;
  wire [63:0] rport_io_ins_331;
  wire [63:0] rport_io_ins_332;
  wire [63:0] rport_io_ins_333;
  wire [63:0] rport_io_ins_334;
  wire [63:0] rport_io_ins_335;
  wire [63:0] rport_io_ins_336;
  wire [63:0] rport_io_ins_337;
  wire [63:0] rport_io_ins_338;
  wire [63:0] rport_io_ins_339;
  wire [63:0] rport_io_ins_340;
  wire [63:0] rport_io_ins_341;
  wire [63:0] rport_io_ins_342;
  wire [63:0] rport_io_ins_343;
  wire [63:0] rport_io_ins_344;
  wire [63:0] rport_io_ins_345;
  wire [63:0] rport_io_ins_346;
  wire [63:0] rport_io_ins_347;
  wire [63:0] rport_io_ins_348;
  wire [63:0] rport_io_ins_349;
  wire [63:0] rport_io_ins_350;
  wire [63:0] rport_io_ins_351;
  wire [63:0] rport_io_ins_352;
  wire [63:0] rport_io_ins_353;
  wire [63:0] rport_io_ins_354;
  wire [63:0] rport_io_ins_355;
  wire [63:0] rport_io_ins_356;
  wire [63:0] rport_io_ins_357;
  wire [63:0] rport_io_ins_358;
  wire [63:0] rport_io_ins_359;
  wire [63:0] rport_io_ins_360;
  wire [63:0] rport_io_ins_361;
  wire [63:0] rport_io_ins_362;
  wire [63:0] rport_io_ins_363;
  wire [63:0] rport_io_ins_364;
  wire [63:0] rport_io_ins_365;
  wire [63:0] rport_io_ins_366;
  wire [63:0] rport_io_ins_367;
  wire [63:0] rport_io_ins_368;
  wire [63:0] rport_io_ins_369;
  wire [63:0] rport_io_ins_370;
  wire [63:0] rport_io_ins_371;
  wire [63:0] rport_io_ins_372;
  wire [63:0] rport_io_ins_373;
  wire [63:0] rport_io_ins_374;
  wire [63:0] rport_io_ins_375;
  wire [63:0] rport_io_ins_376;
  wire [63:0] rport_io_ins_377;
  wire [63:0] rport_io_ins_378;
  wire [63:0] rport_io_ins_379;
  wire [63:0] rport_io_ins_380;
  wire [63:0] rport_io_ins_381;
  wire [63:0] rport_io_ins_382;
  wire [63:0] rport_io_ins_383;
  wire [63:0] rport_io_ins_384;
  wire [63:0] rport_io_ins_385;
  wire [63:0] rport_io_ins_386;
  wire [63:0] rport_io_ins_387;
  wire [63:0] rport_io_ins_388;
  wire [63:0] rport_io_ins_389;
  wire [63:0] rport_io_ins_390;
  wire [63:0] rport_io_ins_391;
  wire [63:0] rport_io_ins_392;
  wire [63:0] rport_io_ins_393;
  wire [63:0] rport_io_ins_394;
  wire [63:0] rport_io_ins_395;
  wire [63:0] rport_io_ins_396;
  wire [63:0] rport_io_ins_397;
  wire [63:0] rport_io_ins_398;
  wire [63:0] rport_io_ins_399;
  wire [63:0] rport_io_ins_400;
  wire [63:0] rport_io_ins_401;
  wire [63:0] rport_io_ins_402;
  wire [63:0] rport_io_ins_403;
  wire [63:0] rport_io_ins_404;
  wire [63:0] rport_io_ins_405;
  wire [63:0] rport_io_ins_406;
  wire [63:0] rport_io_ins_407;
  wire [63:0] rport_io_ins_408;
  wire [63:0] rport_io_ins_409;
  wire [63:0] rport_io_ins_410;
  wire [63:0] rport_io_ins_411;
  wire [63:0] rport_io_ins_412;
  wire [63:0] rport_io_ins_413;
  wire [63:0] rport_io_ins_414;
  wire [63:0] rport_io_ins_415;
  wire [63:0] rport_io_ins_416;
  wire [63:0] rport_io_ins_417;
  wire [63:0] rport_io_ins_418;
  wire [63:0] rport_io_ins_419;
  wire [63:0] rport_io_ins_420;
  wire [63:0] rport_io_ins_421;
  wire [63:0] rport_io_ins_422;
  wire [63:0] rport_io_ins_423;
  wire [63:0] rport_io_ins_424;
  wire [63:0] rport_io_ins_425;
  wire [63:0] rport_io_ins_426;
  wire [63:0] rport_io_ins_427;
  wire [63:0] rport_io_ins_428;
  wire [63:0] rport_io_ins_429;
  wire [63:0] rport_io_ins_430;
  wire [63:0] rport_io_ins_431;
  wire [63:0] rport_io_ins_432;
  wire [63:0] rport_io_ins_433;
  wire [63:0] rport_io_ins_434;
  wire [63:0] rport_io_ins_435;
  wire [63:0] rport_io_ins_436;
  wire [63:0] rport_io_ins_437;
  wire [63:0] rport_io_ins_438;
  wire [63:0] rport_io_ins_439;
  wire [63:0] rport_io_ins_440;
  wire [63:0] rport_io_ins_441;
  wire [63:0] rport_io_ins_442;
  wire [63:0] rport_io_ins_443;
  wire [63:0] rport_io_ins_444;
  wire [63:0] rport_io_ins_445;
  wire [63:0] rport_io_ins_446;
  wire [63:0] rport_io_ins_447;
  wire [63:0] rport_io_ins_448;
  wire [63:0] rport_io_ins_449;
  wire [63:0] rport_io_ins_450;
  wire [63:0] rport_io_ins_451;
  wire [63:0] rport_io_ins_452;
  wire [63:0] rport_io_ins_453;
  wire [63:0] rport_io_ins_454;
  wire [63:0] rport_io_ins_455;
  wire [63:0] rport_io_ins_456;
  wire [63:0] rport_io_ins_457;
  wire [63:0] rport_io_ins_458;
  wire [63:0] rport_io_ins_459;
  wire [63:0] rport_io_ins_460;
  wire [63:0] rport_io_ins_461;
  wire [63:0] rport_io_ins_462;
  wire [63:0] rport_io_ins_463;
  wire [63:0] rport_io_ins_464;
  wire [63:0] rport_io_ins_465;
  wire [63:0] rport_io_ins_466;
  wire [63:0] rport_io_ins_467;
  wire [63:0] rport_io_ins_468;
  wire [63:0] rport_io_ins_469;
  wire [63:0] rport_io_ins_470;
  wire [63:0] rport_io_ins_471;
  wire [63:0] rport_io_ins_472;
  wire [63:0] rport_io_ins_473;
  wire [63:0] rport_io_ins_474;
  wire [63:0] rport_io_ins_475;
  wire [63:0] rport_io_ins_476;
  wire [63:0] rport_io_ins_477;
  wire [63:0] rport_io_ins_478;
  wire [63:0] rport_io_ins_479;
  wire [63:0] rport_io_ins_480;
  wire [63:0] rport_io_ins_481;
  wire [63:0] rport_io_ins_482;
  wire [63:0] rport_io_ins_483;
  wire [63:0] rport_io_ins_484;
  wire [63:0] rport_io_ins_485;
  wire [63:0] rport_io_ins_486;
  wire [63:0] rport_io_ins_487;
  wire [63:0] rport_io_ins_488;
  wire [63:0] rport_io_ins_489;
  wire [63:0] rport_io_ins_490;
  wire [63:0] rport_io_ins_491;
  wire [63:0] rport_io_ins_492;
  wire [63:0] rport_io_ins_493;
  wire [63:0] rport_io_ins_494;
  wire [63:0] rport_io_ins_495;
  wire [63:0] rport_io_ins_496;
  wire [63:0] rport_io_ins_497;
  wire [63:0] rport_io_ins_498;
  wire [63:0] rport_io_ins_499;
  wire [63:0] rport_io_ins_500;
  wire [63:0] rport_io_ins_501;
  wire [63:0] rport_io_ins_502;
  wire [63:0] rport_io_ins_503;
  wire [63:0] rport_io_ins_504;
  wire [63:0] rport_io_ins_505;
  wire [8:0] rport_io_sel;
  wire [63:0] rport_io_out;
  wire [63:0] regOuts_0;
  wire [63:0] regOuts_1;
  wire [63:0] regOuts_2;
  wire [63:0] regOuts_3;
  wire [63:0] regOuts_4;
  wire [63:0] regOuts_5;
  wire [63:0] regOuts_6;
  wire [63:0] regOuts_7;
  wire [63:0] regOuts_8;
  wire [63:0] regOuts_9;
  wire [63:0] regOuts_10;
  wire [63:0] regOuts_11;
  wire [63:0] regOuts_12;
  wire [63:0] regOuts_13;
  wire [63:0] regOuts_14;
  wire [63:0] regOuts_15;
  wire [63:0] regOuts_16;
  wire [63:0] regOuts_17;
  wire [63:0] regOuts_18;
  wire [63:0] regOuts_19;
  wire [63:0] regOuts_20;
  wire [63:0] regOuts_21;
  wire [63:0] regOuts_22;
  wire [63:0] regOuts_23;
  wire [63:0] regOuts_24;
  wire [63:0] regOuts_25;
  wire [63:0] regOuts_26;
  wire [63:0] regOuts_27;
  wire [63:0] regOuts_28;
  wire [63:0] regOuts_29;
  wire [63:0] regOuts_30;
  wire [63:0] regOuts_31;
  wire [63:0] regOuts_32;
  wire [63:0] regOuts_33;
  wire [63:0] regOuts_34;
  wire [63:0] regOuts_35;
  wire [63:0] regOuts_36;
  wire [63:0] regOuts_37;
  wire [63:0] regOuts_38;
  wire [63:0] regOuts_39;
  wire [63:0] regOuts_40;
  wire [63:0] regOuts_41;
  wire [63:0] regOuts_42;
  wire [63:0] regOuts_43;
  wire [63:0] regOuts_44;
  wire [63:0] regOuts_45;
  wire [63:0] regOuts_46;
  wire [63:0] regOuts_47;
  wire [63:0] regOuts_48;
  wire [63:0] regOuts_49;
  wire [63:0] regOuts_50;
  wire [63:0] regOuts_51;
  wire [63:0] regOuts_52;
  wire [63:0] regOuts_53;
  wire [63:0] regOuts_54;
  wire [63:0] regOuts_55;
  wire [63:0] regOuts_56;
  wire [63:0] regOuts_57;
  wire [63:0] regOuts_58;
  wire [63:0] regOuts_59;
  wire [63:0] regOuts_60;
  wire [63:0] regOuts_61;
  wire [63:0] regOuts_62;
  wire [63:0] regOuts_63;
  wire [63:0] regOuts_64;
  wire [63:0] regOuts_65;
  wire [63:0] regOuts_66;
  wire [63:0] regOuts_67;
  wire [63:0] regOuts_68;
  wire [63:0] regOuts_69;
  wire [63:0] regOuts_70;
  wire [63:0] regOuts_71;
  wire [63:0] regOuts_72;
  wire [63:0] regOuts_73;
  wire [63:0] regOuts_74;
  wire [63:0] regOuts_75;
  wire [63:0] regOuts_76;
  wire [63:0] regOuts_77;
  wire [63:0] regOuts_78;
  wire [63:0] regOuts_79;
  wire [63:0] regOuts_80;
  wire [63:0] regOuts_81;
  wire [63:0] regOuts_82;
  wire [63:0] regOuts_83;
  wire [63:0] regOuts_84;
  wire [63:0] regOuts_85;
  wire [63:0] regOuts_86;
  wire [63:0] regOuts_87;
  wire [63:0] regOuts_88;
  wire [63:0] regOuts_89;
  wire [63:0] regOuts_90;
  wire [63:0] regOuts_91;
  wire [63:0] regOuts_92;
  wire [63:0] regOuts_93;
  wire [63:0] regOuts_94;
  wire [63:0] regOuts_95;
  wire [63:0] regOuts_96;
  wire [63:0] regOuts_97;
  wire [63:0] regOuts_98;
  wire [63:0] regOuts_99;
  wire [63:0] regOuts_100;
  wire [63:0] regOuts_101;
  wire [63:0] regOuts_102;
  wire [63:0] regOuts_103;
  wire [63:0] regOuts_104;
  wire [63:0] regOuts_105;
  wire [63:0] regOuts_106;
  wire [63:0] regOuts_107;
  wire [63:0] regOuts_108;
  wire [63:0] regOuts_109;
  wire [63:0] regOuts_110;
  wire [63:0] regOuts_111;
  wire [63:0] regOuts_112;
  wire [63:0] regOuts_113;
  wire [63:0] regOuts_114;
  wire [63:0] regOuts_115;
  wire [63:0] regOuts_116;
  wire [63:0] regOuts_117;
  wire [63:0] regOuts_118;
  wire [63:0] regOuts_119;
  wire [63:0] regOuts_120;
  wire [63:0] regOuts_121;
  wire [63:0] regOuts_122;
  wire [63:0] regOuts_123;
  wire [63:0] regOuts_124;
  wire [63:0] regOuts_125;
  wire [63:0] regOuts_126;
  wire [63:0] regOuts_127;
  wire [63:0] regOuts_128;
  wire [63:0] regOuts_129;
  wire [63:0] regOuts_130;
  wire [63:0] regOuts_131;
  wire [63:0] regOuts_132;
  wire [63:0] regOuts_133;
  wire [63:0] regOuts_134;
  wire [63:0] regOuts_135;
  wire [63:0] regOuts_136;
  wire [63:0] regOuts_137;
  wire [63:0] regOuts_138;
  wire [63:0] regOuts_139;
  wire [63:0] regOuts_140;
  wire [63:0] regOuts_141;
  wire [63:0] regOuts_142;
  wire [63:0] regOuts_143;
  wire [63:0] regOuts_144;
  wire [63:0] regOuts_145;
  wire [63:0] regOuts_146;
  wire [63:0] regOuts_147;
  wire [63:0] regOuts_148;
  wire [63:0] regOuts_149;
  wire [63:0] regOuts_150;
  wire [63:0] regOuts_151;
  wire [63:0] regOuts_152;
  wire [63:0] regOuts_153;
  wire [63:0] regOuts_154;
  wire [63:0] regOuts_155;
  wire [63:0] regOuts_156;
  wire [63:0] regOuts_157;
  wire [63:0] regOuts_158;
  wire [63:0] regOuts_159;
  wire [63:0] regOuts_160;
  wire [63:0] regOuts_161;
  wire [63:0] regOuts_162;
  wire [63:0] regOuts_163;
  wire [63:0] regOuts_164;
  wire [63:0] regOuts_165;
  wire [63:0] regOuts_166;
  wire [63:0] regOuts_167;
  wire [63:0] regOuts_168;
  wire [63:0] regOuts_169;
  wire [63:0] regOuts_170;
  wire [63:0] regOuts_171;
  wire [63:0] regOuts_172;
  wire [63:0] regOuts_173;
  wire [63:0] regOuts_174;
  wire [63:0] regOuts_175;
  wire [63:0] regOuts_176;
  wire [63:0] regOuts_177;
  wire [63:0] regOuts_178;
  wire [63:0] regOuts_179;
  wire [63:0] regOuts_180;
  wire [63:0] regOuts_181;
  wire [63:0] regOuts_182;
  wire [63:0] regOuts_183;
  wire [63:0] regOuts_184;
  wire [63:0] regOuts_185;
  wire [63:0] regOuts_186;
  wire [63:0] regOuts_187;
  wire [63:0] regOuts_188;
  wire [63:0] regOuts_189;
  wire [63:0] regOuts_190;
  wire [63:0] regOuts_191;
  wire [63:0] regOuts_192;
  wire [63:0] regOuts_193;
  wire [63:0] regOuts_194;
  wire [63:0] regOuts_195;
  wire [63:0] regOuts_196;
  wire [63:0] regOuts_197;
  wire [63:0] regOuts_198;
  wire [63:0] regOuts_199;
  wire [63:0] regOuts_200;
  wire [63:0] regOuts_201;
  wire [63:0] regOuts_202;
  wire [63:0] regOuts_203;
  wire [63:0] regOuts_204;
  wire [63:0] regOuts_205;
  wire [63:0] regOuts_206;
  wire [63:0] regOuts_207;
  wire [63:0] regOuts_208;
  wire [63:0] regOuts_209;
  wire [63:0] regOuts_210;
  wire [63:0] regOuts_211;
  wire [63:0] regOuts_212;
  wire [63:0] regOuts_213;
  wire [63:0] regOuts_214;
  wire [63:0] regOuts_215;
  wire [63:0] regOuts_216;
  wire [63:0] regOuts_217;
  wire [63:0] regOuts_218;
  wire [63:0] regOuts_219;
  wire [63:0] regOuts_220;
  wire [63:0] regOuts_221;
  wire [63:0] regOuts_222;
  wire [63:0] regOuts_223;
  wire [63:0] regOuts_224;
  wire [63:0] regOuts_225;
  wire [63:0] regOuts_226;
  wire [63:0] regOuts_227;
  wire [63:0] regOuts_228;
  wire [63:0] regOuts_229;
  wire [63:0] regOuts_230;
  wire [63:0] regOuts_231;
  wire [63:0] regOuts_232;
  wire [63:0] regOuts_233;
  wire [63:0] regOuts_234;
  wire [63:0] regOuts_235;
  wire [63:0] regOuts_236;
  wire [63:0] regOuts_237;
  wire [63:0] regOuts_238;
  wire [63:0] regOuts_239;
  wire [63:0] regOuts_240;
  wire [63:0] regOuts_241;
  wire [63:0] regOuts_242;
  wire [63:0] regOuts_243;
  wire [63:0] regOuts_244;
  wire [63:0] regOuts_245;
  wire [63:0] regOuts_246;
  wire [63:0] regOuts_247;
  wire [63:0] regOuts_248;
  wire [63:0] regOuts_249;
  wire [63:0] regOuts_250;
  wire [63:0] regOuts_251;
  wire [63:0] regOuts_252;
  wire [63:0] regOuts_253;
  wire [63:0] regOuts_254;
  wire [63:0] regOuts_255;
  wire [63:0] regOuts_256;
  wire [63:0] regOuts_257;
  wire [63:0] regOuts_258;
  wire [63:0] regOuts_259;
  wire [63:0] regOuts_260;
  wire [63:0] regOuts_261;
  wire [63:0] regOuts_262;
  wire [63:0] regOuts_263;
  wire [63:0] regOuts_264;
  wire [63:0] regOuts_265;
  wire [63:0] regOuts_266;
  wire [63:0] regOuts_267;
  wire [63:0] regOuts_268;
  wire [63:0] regOuts_269;
  wire [63:0] regOuts_270;
  wire [63:0] regOuts_271;
  wire [63:0] regOuts_272;
  wire [63:0] regOuts_273;
  wire [63:0] regOuts_274;
  wire [63:0] regOuts_275;
  wire [63:0] regOuts_276;
  wire [63:0] regOuts_277;
  wire [63:0] regOuts_278;
  wire [63:0] regOuts_279;
  wire [63:0] regOuts_280;
  wire [63:0] regOuts_281;
  wire [63:0] regOuts_282;
  wire [63:0] regOuts_283;
  wire [63:0] regOuts_284;
  wire [63:0] regOuts_285;
  wire [63:0] regOuts_286;
  wire [63:0] regOuts_287;
  wire [63:0] regOuts_288;
  wire [63:0] regOuts_289;
  wire [63:0] regOuts_290;
  wire [63:0] regOuts_291;
  wire [63:0] regOuts_292;
  wire [63:0] regOuts_293;
  wire [63:0] regOuts_294;
  wire [63:0] regOuts_295;
  wire [63:0] regOuts_296;
  wire [63:0] regOuts_297;
  wire [63:0] regOuts_298;
  wire [63:0] regOuts_299;
  wire [63:0] regOuts_300;
  wire [63:0] regOuts_301;
  wire [63:0] regOuts_302;
  wire [63:0] regOuts_303;
  wire [63:0] regOuts_304;
  wire [63:0] regOuts_305;
  wire [63:0] regOuts_306;
  wire [63:0] regOuts_307;
  wire [63:0] regOuts_308;
  wire [63:0] regOuts_309;
  wire [63:0] regOuts_310;
  wire [63:0] regOuts_311;
  wire [63:0] regOuts_312;
  wire [63:0] regOuts_313;
  wire [63:0] regOuts_314;
  wire [63:0] regOuts_315;
  wire [63:0] regOuts_316;
  wire [63:0] regOuts_317;
  wire [63:0] regOuts_318;
  wire [63:0] regOuts_319;
  wire [63:0] regOuts_320;
  wire [63:0] regOuts_321;
  wire [63:0] regOuts_322;
  wire [63:0] regOuts_323;
  wire [63:0] regOuts_324;
  wire [63:0] regOuts_325;
  wire [63:0] regOuts_326;
  wire [63:0] regOuts_327;
  wire [63:0] regOuts_328;
  wire [63:0] regOuts_329;
  wire [63:0] regOuts_330;
  wire [63:0] regOuts_331;
  wire [63:0] regOuts_332;
  wire [63:0] regOuts_333;
  wire [63:0] regOuts_334;
  wire [63:0] regOuts_335;
  wire [63:0] regOuts_336;
  wire [63:0] regOuts_337;
  wire [63:0] regOuts_338;
  wire [63:0] regOuts_339;
  wire [63:0] regOuts_340;
  wire [63:0] regOuts_341;
  wire [63:0] regOuts_342;
  wire [63:0] regOuts_343;
  wire [63:0] regOuts_344;
  wire [63:0] regOuts_345;
  wire [63:0] regOuts_346;
  wire [63:0] regOuts_347;
  wire [63:0] regOuts_348;
  wire [63:0] regOuts_349;
  wire [63:0] regOuts_350;
  wire [63:0] regOuts_351;
  wire [63:0] regOuts_352;
  wire [63:0] regOuts_353;
  wire [63:0] regOuts_354;
  wire [63:0] regOuts_355;
  wire [63:0] regOuts_356;
  wire [63:0] regOuts_357;
  wire [63:0] regOuts_358;
  wire [63:0] regOuts_359;
  wire [63:0] regOuts_360;
  wire [63:0] regOuts_361;
  wire [63:0] regOuts_362;
  wire [63:0] regOuts_363;
  wire [63:0] regOuts_364;
  wire [63:0] regOuts_365;
  wire [63:0] regOuts_366;
  wire [63:0] regOuts_367;
  wire [63:0] regOuts_368;
  wire [63:0] regOuts_369;
  wire [63:0] regOuts_370;
  wire [63:0] regOuts_371;
  wire [63:0] regOuts_372;
  wire [63:0] regOuts_373;
  wire [63:0] regOuts_374;
  wire [63:0] regOuts_375;
  wire [63:0] regOuts_376;
  wire [63:0] regOuts_377;
  wire [63:0] regOuts_378;
  wire [63:0] regOuts_379;
  wire [63:0] regOuts_380;
  wire [63:0] regOuts_381;
  wire [63:0] regOuts_382;
  wire [63:0] regOuts_383;
  wire [63:0] regOuts_384;
  wire [63:0] regOuts_385;
  wire [63:0] regOuts_386;
  wire [63:0] regOuts_387;
  wire [63:0] regOuts_388;
  wire [63:0] regOuts_389;
  wire [63:0] regOuts_390;
  wire [63:0] regOuts_391;
  wire [63:0] regOuts_392;
  wire [63:0] regOuts_393;
  wire [63:0] regOuts_394;
  wire [63:0] regOuts_395;
  wire [63:0] regOuts_396;
  wire [63:0] regOuts_397;
  wire [63:0] regOuts_398;
  wire [63:0] regOuts_399;
  wire [63:0] regOuts_400;
  wire [63:0] regOuts_401;
  wire [63:0] regOuts_402;
  wire [63:0] regOuts_403;
  wire [63:0] regOuts_404;
  wire [63:0] regOuts_405;
  wire [63:0] regOuts_406;
  wire [63:0] regOuts_407;
  wire [63:0] regOuts_408;
  wire [63:0] regOuts_409;
  wire [63:0] regOuts_410;
  wire [63:0] regOuts_411;
  wire [63:0] regOuts_412;
  wire [63:0] regOuts_413;
  wire [63:0] regOuts_414;
  wire [63:0] regOuts_415;
  wire [63:0] regOuts_416;
  wire [63:0] regOuts_417;
  wire [63:0] regOuts_418;
  wire [63:0] regOuts_419;
  wire [63:0] regOuts_420;
  wire [63:0] regOuts_421;
  wire [63:0] regOuts_422;
  wire [63:0] regOuts_423;
  wire [63:0] regOuts_424;
  wire [63:0] regOuts_425;
  wire [63:0] regOuts_426;
  wire [63:0] regOuts_427;
  wire [63:0] regOuts_428;
  wire [63:0] regOuts_429;
  wire [63:0] regOuts_430;
  wire [63:0] regOuts_431;
  wire [63:0] regOuts_432;
  wire [63:0] regOuts_433;
  wire [63:0] regOuts_434;
  wire [63:0] regOuts_435;
  wire [63:0] regOuts_436;
  wire [63:0] regOuts_437;
  wire [63:0] regOuts_438;
  wire [63:0] regOuts_439;
  wire [63:0] regOuts_440;
  wire [63:0] regOuts_441;
  wire [63:0] regOuts_442;
  wire [63:0] regOuts_443;
  wire [63:0] regOuts_444;
  wire [63:0] regOuts_445;
  wire [63:0] regOuts_446;
  wire [63:0] regOuts_447;
  wire [63:0] regOuts_448;
  wire [63:0] regOuts_449;
  wire [63:0] regOuts_450;
  wire [63:0] regOuts_451;
  wire [63:0] regOuts_452;
  wire [63:0] regOuts_453;
  wire [63:0] regOuts_454;
  wire [63:0] regOuts_455;
  wire [63:0] regOuts_456;
  wire [63:0] regOuts_457;
  wire [63:0] regOuts_458;
  wire [63:0] regOuts_459;
  wire [63:0] regOuts_460;
  wire [63:0] regOuts_461;
  wire [63:0] regOuts_462;
  wire [63:0] regOuts_463;
  wire [63:0] regOuts_464;
  wire [63:0] regOuts_465;
  wire [63:0] regOuts_466;
  wire [63:0] regOuts_467;
  wire [63:0] regOuts_468;
  wire [63:0] regOuts_469;
  wire [63:0] regOuts_470;
  wire [63:0] regOuts_471;
  wire [63:0] regOuts_472;
  wire [63:0] regOuts_473;
  wire [63:0] regOuts_474;
  wire [63:0] regOuts_475;
  wire [63:0] regOuts_476;
  wire [63:0] regOuts_477;
  wire [63:0] regOuts_478;
  wire [63:0] regOuts_479;
  wire [63:0] regOuts_480;
  wire [63:0] regOuts_481;
  wire [63:0] regOuts_482;
  wire [63:0] regOuts_483;
  wire [63:0] regOuts_484;
  wire [63:0] regOuts_485;
  wire [63:0] regOuts_486;
  wire [63:0] regOuts_487;
  wire [63:0] regOuts_488;
  wire [63:0] regOuts_489;
  wire [63:0] regOuts_490;
  wire [63:0] regOuts_491;
  wire [63:0] regOuts_492;
  wire [63:0] regOuts_493;
  wire [63:0] regOuts_494;
  wire [63:0] regOuts_495;
  wire [63:0] regOuts_496;
  wire [63:0] regOuts_497;
  wire [63:0] regOuts_498;
  wire [63:0] regOuts_499;
  wire [63:0] regOuts_500;
  wire [63:0] regOuts_501;
  wire [63:0] regOuts_502;
  wire [63:0] regOuts_503;
  wire [63:0] regOuts_504;
  wire [63:0] regOuts_505;
  wire [31:0] _T_5611;
  wire  _T_5612;
  wire [31:0] _T_5613;
  wire [31:0] _T_5614;
  wire [31:0] _T_5615;
  wire [63:0] _T_5618_0;
  wire [63:0] _T_5618_1;
  wire [63:0] _T_5618_2;
  wire [63:0] _T_5618_3;
  wire [63:0] _T_5618_4;
  FF_136 regs_0 (
    .clock(regs_0_clock),
    .reset(regs_0_reset),
    .io_in(regs_0_io_in),
    .io_init(regs_0_io_init),
    .io_reset(regs_0_io_reset),
    .io_out(regs_0_io_out),
    .io_enable(regs_0_io_enable)
  );
  FF_136 regs_1 (
    .clock(regs_1_clock),
    .reset(regs_1_reset),
    .io_in(regs_1_io_in),
    .io_init(regs_1_io_init),
    .io_reset(regs_1_io_reset),
    .io_out(regs_1_io_out),
    .io_enable(regs_1_io_enable)
  );
  FF_136 regs_2 (
    .clock(regs_2_clock),
    .reset(regs_2_reset),
    .io_in(regs_2_io_in),
    .io_init(regs_2_io_init),
    .io_reset(regs_2_io_reset),
    .io_out(regs_2_io_out),
    .io_enable(regs_2_io_enable)
  );
  FF_136 regs_3 (
    .clock(regs_3_clock),
    .reset(regs_3_reset),
    .io_in(regs_3_io_in),
    .io_init(regs_3_io_init),
    .io_reset(regs_3_io_reset),
    .io_out(regs_3_io_out),
    .io_enable(regs_3_io_enable)
  );
  FF_136 regs_4 (
    .clock(regs_4_clock),
    .reset(regs_4_reset),
    .io_in(regs_4_io_in),
    .io_init(regs_4_io_init),
    .io_reset(regs_4_io_reset),
    .io_out(regs_4_io_out),
    .io_enable(regs_4_io_enable)
  );
  FF_136 regs_5 (
    .clock(regs_5_clock),
    .reset(regs_5_reset),
    .io_in(regs_5_io_in),
    .io_init(regs_5_io_init),
    .io_reset(regs_5_io_reset),
    .io_out(regs_5_io_out),
    .io_enable(regs_5_io_enable)
  );
  FF_136 regs_6 (
    .clock(regs_6_clock),
    .reset(regs_6_reset),
    .io_in(regs_6_io_in),
    .io_init(regs_6_io_init),
    .io_reset(regs_6_io_reset),
    .io_out(regs_6_io_out),
    .io_enable(regs_6_io_enable)
  );
  FF_136 regs_7 (
    .clock(regs_7_clock),
    .reset(regs_7_reset),
    .io_in(regs_7_io_in),
    .io_init(regs_7_io_init),
    .io_reset(regs_7_io_reset),
    .io_out(regs_7_io_out),
    .io_enable(regs_7_io_enable)
  );
  FF_136 regs_8 (
    .clock(regs_8_clock),
    .reset(regs_8_reset),
    .io_in(regs_8_io_in),
    .io_init(regs_8_io_init),
    .io_reset(regs_8_io_reset),
    .io_out(regs_8_io_out),
    .io_enable(regs_8_io_enable)
  );
  FF_136 regs_9 (
    .clock(regs_9_clock),
    .reset(regs_9_reset),
    .io_in(regs_9_io_in),
    .io_init(regs_9_io_init),
    .io_reset(regs_9_io_reset),
    .io_out(regs_9_io_out),
    .io_enable(regs_9_io_enable)
  );
  FF_136 regs_10 (
    .clock(regs_10_clock),
    .reset(regs_10_reset),
    .io_in(regs_10_io_in),
    .io_init(regs_10_io_init),
    .io_reset(regs_10_io_reset),
    .io_out(regs_10_io_out),
    .io_enable(regs_10_io_enable)
  );
  FF_136 regs_11 (
    .clock(regs_11_clock),
    .reset(regs_11_reset),
    .io_in(regs_11_io_in),
    .io_init(regs_11_io_init),
    .io_reset(regs_11_io_reset),
    .io_out(regs_11_io_out),
    .io_enable(regs_11_io_enable)
  );
  FF_136 regs_12 (
    .clock(regs_12_clock),
    .reset(regs_12_reset),
    .io_in(regs_12_io_in),
    .io_init(regs_12_io_init),
    .io_reset(regs_12_io_reset),
    .io_out(regs_12_io_out),
    .io_enable(regs_12_io_enable)
  );
  FF_136 regs_13 (
    .clock(regs_13_clock),
    .reset(regs_13_reset),
    .io_in(regs_13_io_in),
    .io_init(regs_13_io_init),
    .io_reset(regs_13_io_reset),
    .io_out(regs_13_io_out),
    .io_enable(regs_13_io_enable)
  );
  FF_136 regs_14 (
    .clock(regs_14_clock),
    .reset(regs_14_reset),
    .io_in(regs_14_io_in),
    .io_init(regs_14_io_init),
    .io_reset(regs_14_io_reset),
    .io_out(regs_14_io_out),
    .io_enable(regs_14_io_enable)
  );
  FF_136 regs_15 (
    .clock(regs_15_clock),
    .reset(regs_15_reset),
    .io_in(regs_15_io_in),
    .io_init(regs_15_io_init),
    .io_reset(regs_15_io_reset),
    .io_out(regs_15_io_out),
    .io_enable(regs_15_io_enable)
  );
  FF_136 regs_16 (
    .clock(regs_16_clock),
    .reset(regs_16_reset),
    .io_in(regs_16_io_in),
    .io_init(regs_16_io_init),
    .io_reset(regs_16_io_reset),
    .io_out(regs_16_io_out),
    .io_enable(regs_16_io_enable)
  );
  FF_136 regs_17 (
    .clock(regs_17_clock),
    .reset(regs_17_reset),
    .io_in(regs_17_io_in),
    .io_init(regs_17_io_init),
    .io_reset(regs_17_io_reset),
    .io_out(regs_17_io_out),
    .io_enable(regs_17_io_enable)
  );
  FF_136 regs_18 (
    .clock(regs_18_clock),
    .reset(regs_18_reset),
    .io_in(regs_18_io_in),
    .io_init(regs_18_io_init),
    .io_reset(regs_18_io_reset),
    .io_out(regs_18_io_out),
    .io_enable(regs_18_io_enable)
  );
  FF_136 regs_19 (
    .clock(regs_19_clock),
    .reset(regs_19_reset),
    .io_in(regs_19_io_in),
    .io_init(regs_19_io_init),
    .io_reset(regs_19_io_reset),
    .io_out(regs_19_io_out),
    .io_enable(regs_19_io_enable)
  );
  FF_136 regs_20 (
    .clock(regs_20_clock),
    .reset(regs_20_reset),
    .io_in(regs_20_io_in),
    .io_init(regs_20_io_init),
    .io_reset(regs_20_io_reset),
    .io_out(regs_20_io_out),
    .io_enable(regs_20_io_enable)
  );
  FF_136 regs_21 (
    .clock(regs_21_clock),
    .reset(regs_21_reset),
    .io_in(regs_21_io_in),
    .io_init(regs_21_io_init),
    .io_reset(regs_21_io_reset),
    .io_out(regs_21_io_out),
    .io_enable(regs_21_io_enable)
  );
  FF_136 regs_22 (
    .clock(regs_22_clock),
    .reset(regs_22_reset),
    .io_in(regs_22_io_in),
    .io_init(regs_22_io_init),
    .io_reset(regs_22_io_reset),
    .io_out(regs_22_io_out),
    .io_enable(regs_22_io_enable)
  );
  FF_136 regs_23 (
    .clock(regs_23_clock),
    .reset(regs_23_reset),
    .io_in(regs_23_io_in),
    .io_init(regs_23_io_init),
    .io_reset(regs_23_io_reset),
    .io_out(regs_23_io_out),
    .io_enable(regs_23_io_enable)
  );
  FF_136 regs_24 (
    .clock(regs_24_clock),
    .reset(regs_24_reset),
    .io_in(regs_24_io_in),
    .io_init(regs_24_io_init),
    .io_reset(regs_24_io_reset),
    .io_out(regs_24_io_out),
    .io_enable(regs_24_io_enable)
  );
  FF_136 regs_25 (
    .clock(regs_25_clock),
    .reset(regs_25_reset),
    .io_in(regs_25_io_in),
    .io_init(regs_25_io_init),
    .io_reset(regs_25_io_reset),
    .io_out(regs_25_io_out),
    .io_enable(regs_25_io_enable)
  );
  FF_136 regs_26 (
    .clock(regs_26_clock),
    .reset(regs_26_reset),
    .io_in(regs_26_io_in),
    .io_init(regs_26_io_init),
    .io_reset(regs_26_io_reset),
    .io_out(regs_26_io_out),
    .io_enable(regs_26_io_enable)
  );
  FF_136 regs_27 (
    .clock(regs_27_clock),
    .reset(regs_27_reset),
    .io_in(regs_27_io_in),
    .io_init(regs_27_io_init),
    .io_reset(regs_27_io_reset),
    .io_out(regs_27_io_out),
    .io_enable(regs_27_io_enable)
  );
  FF_136 regs_28 (
    .clock(regs_28_clock),
    .reset(regs_28_reset),
    .io_in(regs_28_io_in),
    .io_init(regs_28_io_init),
    .io_reset(regs_28_io_reset),
    .io_out(regs_28_io_out),
    .io_enable(regs_28_io_enable)
  );
  FF_136 regs_29 (
    .clock(regs_29_clock),
    .reset(regs_29_reset),
    .io_in(regs_29_io_in),
    .io_init(regs_29_io_init),
    .io_reset(regs_29_io_reset),
    .io_out(regs_29_io_out),
    .io_enable(regs_29_io_enable)
  );
  FF_136 regs_30 (
    .clock(regs_30_clock),
    .reset(regs_30_reset),
    .io_in(regs_30_io_in),
    .io_init(regs_30_io_init),
    .io_reset(regs_30_io_reset),
    .io_out(regs_30_io_out),
    .io_enable(regs_30_io_enable)
  );
  FF_136 regs_31 (
    .clock(regs_31_clock),
    .reset(regs_31_reset),
    .io_in(regs_31_io_in),
    .io_init(regs_31_io_init),
    .io_reset(regs_31_io_reset),
    .io_out(regs_31_io_out),
    .io_enable(regs_31_io_enable)
  );
  FF_136 regs_32 (
    .clock(regs_32_clock),
    .reset(regs_32_reset),
    .io_in(regs_32_io_in),
    .io_init(regs_32_io_init),
    .io_reset(regs_32_io_reset),
    .io_out(regs_32_io_out),
    .io_enable(regs_32_io_enable)
  );
  FF_136 regs_33 (
    .clock(regs_33_clock),
    .reset(regs_33_reset),
    .io_in(regs_33_io_in),
    .io_init(regs_33_io_init),
    .io_reset(regs_33_io_reset),
    .io_out(regs_33_io_out),
    .io_enable(regs_33_io_enable)
  );
  FF_136 regs_34 (
    .clock(regs_34_clock),
    .reset(regs_34_reset),
    .io_in(regs_34_io_in),
    .io_init(regs_34_io_init),
    .io_reset(regs_34_io_reset),
    .io_out(regs_34_io_out),
    .io_enable(regs_34_io_enable)
  );
  FF_136 regs_35 (
    .clock(regs_35_clock),
    .reset(regs_35_reset),
    .io_in(regs_35_io_in),
    .io_init(regs_35_io_init),
    .io_reset(regs_35_io_reset),
    .io_out(regs_35_io_out),
    .io_enable(regs_35_io_enable)
  );
  FF_136 regs_36 (
    .clock(regs_36_clock),
    .reset(regs_36_reset),
    .io_in(regs_36_io_in),
    .io_init(regs_36_io_init),
    .io_reset(regs_36_io_reset),
    .io_out(regs_36_io_out),
    .io_enable(regs_36_io_enable)
  );
  FF_136 regs_37 (
    .clock(regs_37_clock),
    .reset(regs_37_reset),
    .io_in(regs_37_io_in),
    .io_init(regs_37_io_init),
    .io_reset(regs_37_io_reset),
    .io_out(regs_37_io_out),
    .io_enable(regs_37_io_enable)
  );
  FF_136 regs_38 (
    .clock(regs_38_clock),
    .reset(regs_38_reset),
    .io_in(regs_38_io_in),
    .io_init(regs_38_io_init),
    .io_reset(regs_38_io_reset),
    .io_out(regs_38_io_out),
    .io_enable(regs_38_io_enable)
  );
  FF_136 regs_39 (
    .clock(regs_39_clock),
    .reset(regs_39_reset),
    .io_in(regs_39_io_in),
    .io_init(regs_39_io_init),
    .io_reset(regs_39_io_reset),
    .io_out(regs_39_io_out),
    .io_enable(regs_39_io_enable)
  );
  FF_136 regs_40 (
    .clock(regs_40_clock),
    .reset(regs_40_reset),
    .io_in(regs_40_io_in),
    .io_init(regs_40_io_init),
    .io_reset(regs_40_io_reset),
    .io_out(regs_40_io_out),
    .io_enable(regs_40_io_enable)
  );
  FF_136 regs_41 (
    .clock(regs_41_clock),
    .reset(regs_41_reset),
    .io_in(regs_41_io_in),
    .io_init(regs_41_io_init),
    .io_reset(regs_41_io_reset),
    .io_out(regs_41_io_out),
    .io_enable(regs_41_io_enable)
  );
  FF_136 regs_42 (
    .clock(regs_42_clock),
    .reset(regs_42_reset),
    .io_in(regs_42_io_in),
    .io_init(regs_42_io_init),
    .io_reset(regs_42_io_reset),
    .io_out(regs_42_io_out),
    .io_enable(regs_42_io_enable)
  );
  FF_136 regs_43 (
    .clock(regs_43_clock),
    .reset(regs_43_reset),
    .io_in(regs_43_io_in),
    .io_init(regs_43_io_init),
    .io_reset(regs_43_io_reset),
    .io_out(regs_43_io_out),
    .io_enable(regs_43_io_enable)
  );
  FF_136 regs_44 (
    .clock(regs_44_clock),
    .reset(regs_44_reset),
    .io_in(regs_44_io_in),
    .io_init(regs_44_io_init),
    .io_reset(regs_44_io_reset),
    .io_out(regs_44_io_out),
    .io_enable(regs_44_io_enable)
  );
  FF_136 regs_45 (
    .clock(regs_45_clock),
    .reset(regs_45_reset),
    .io_in(regs_45_io_in),
    .io_init(regs_45_io_init),
    .io_reset(regs_45_io_reset),
    .io_out(regs_45_io_out),
    .io_enable(regs_45_io_enable)
  );
  FF_136 regs_46 (
    .clock(regs_46_clock),
    .reset(regs_46_reset),
    .io_in(regs_46_io_in),
    .io_init(regs_46_io_init),
    .io_reset(regs_46_io_reset),
    .io_out(regs_46_io_out),
    .io_enable(regs_46_io_enable)
  );
  FF_136 regs_47 (
    .clock(regs_47_clock),
    .reset(regs_47_reset),
    .io_in(regs_47_io_in),
    .io_init(regs_47_io_init),
    .io_reset(regs_47_io_reset),
    .io_out(regs_47_io_out),
    .io_enable(regs_47_io_enable)
  );
  FF_136 regs_48 (
    .clock(regs_48_clock),
    .reset(regs_48_reset),
    .io_in(regs_48_io_in),
    .io_init(regs_48_io_init),
    .io_reset(regs_48_io_reset),
    .io_out(regs_48_io_out),
    .io_enable(regs_48_io_enable)
  );
  FF_136 regs_49 (
    .clock(regs_49_clock),
    .reset(regs_49_reset),
    .io_in(regs_49_io_in),
    .io_init(regs_49_io_init),
    .io_reset(regs_49_io_reset),
    .io_out(regs_49_io_out),
    .io_enable(regs_49_io_enable)
  );
  FF_136 regs_50 (
    .clock(regs_50_clock),
    .reset(regs_50_reset),
    .io_in(regs_50_io_in),
    .io_init(regs_50_io_init),
    .io_reset(regs_50_io_reset),
    .io_out(regs_50_io_out),
    .io_enable(regs_50_io_enable)
  );
  FF_136 regs_51 (
    .clock(regs_51_clock),
    .reset(regs_51_reset),
    .io_in(regs_51_io_in),
    .io_init(regs_51_io_init),
    .io_reset(regs_51_io_reset),
    .io_out(regs_51_io_out),
    .io_enable(regs_51_io_enable)
  );
  FF_136 regs_52 (
    .clock(regs_52_clock),
    .reset(regs_52_reset),
    .io_in(regs_52_io_in),
    .io_init(regs_52_io_init),
    .io_reset(regs_52_io_reset),
    .io_out(regs_52_io_out),
    .io_enable(regs_52_io_enable)
  );
  FF_136 regs_53 (
    .clock(regs_53_clock),
    .reset(regs_53_reset),
    .io_in(regs_53_io_in),
    .io_init(regs_53_io_init),
    .io_reset(regs_53_io_reset),
    .io_out(regs_53_io_out),
    .io_enable(regs_53_io_enable)
  );
  FF_136 regs_54 (
    .clock(regs_54_clock),
    .reset(regs_54_reset),
    .io_in(regs_54_io_in),
    .io_init(regs_54_io_init),
    .io_reset(regs_54_io_reset),
    .io_out(regs_54_io_out),
    .io_enable(regs_54_io_enable)
  );
  FF_136 regs_55 (
    .clock(regs_55_clock),
    .reset(regs_55_reset),
    .io_in(regs_55_io_in),
    .io_init(regs_55_io_init),
    .io_reset(regs_55_io_reset),
    .io_out(regs_55_io_out),
    .io_enable(regs_55_io_enable)
  );
  FF_136 regs_56 (
    .clock(regs_56_clock),
    .reset(regs_56_reset),
    .io_in(regs_56_io_in),
    .io_init(regs_56_io_init),
    .io_reset(regs_56_io_reset),
    .io_out(regs_56_io_out),
    .io_enable(regs_56_io_enable)
  );
  FF_136 regs_57 (
    .clock(regs_57_clock),
    .reset(regs_57_reset),
    .io_in(regs_57_io_in),
    .io_init(regs_57_io_init),
    .io_reset(regs_57_io_reset),
    .io_out(regs_57_io_out),
    .io_enable(regs_57_io_enable)
  );
  FF_136 regs_58 (
    .clock(regs_58_clock),
    .reset(regs_58_reset),
    .io_in(regs_58_io_in),
    .io_init(regs_58_io_init),
    .io_reset(regs_58_io_reset),
    .io_out(regs_58_io_out),
    .io_enable(regs_58_io_enable)
  );
  FF_136 regs_59 (
    .clock(regs_59_clock),
    .reset(regs_59_reset),
    .io_in(regs_59_io_in),
    .io_init(regs_59_io_init),
    .io_reset(regs_59_io_reset),
    .io_out(regs_59_io_out),
    .io_enable(regs_59_io_enable)
  );
  FF_136 regs_60 (
    .clock(regs_60_clock),
    .reset(regs_60_reset),
    .io_in(regs_60_io_in),
    .io_init(regs_60_io_init),
    .io_reset(regs_60_io_reset),
    .io_out(regs_60_io_out),
    .io_enable(regs_60_io_enable)
  );
  FF_136 regs_61 (
    .clock(regs_61_clock),
    .reset(regs_61_reset),
    .io_in(regs_61_io_in),
    .io_init(regs_61_io_init),
    .io_reset(regs_61_io_reset),
    .io_out(regs_61_io_out),
    .io_enable(regs_61_io_enable)
  );
  FF_136 regs_62 (
    .clock(regs_62_clock),
    .reset(regs_62_reset),
    .io_in(regs_62_io_in),
    .io_init(regs_62_io_init),
    .io_reset(regs_62_io_reset),
    .io_out(regs_62_io_out),
    .io_enable(regs_62_io_enable)
  );
  FF_136 regs_63 (
    .clock(regs_63_clock),
    .reset(regs_63_reset),
    .io_in(regs_63_io_in),
    .io_init(regs_63_io_init),
    .io_reset(regs_63_io_reset),
    .io_out(regs_63_io_out),
    .io_enable(regs_63_io_enable)
  );
  FF_136 regs_64 (
    .clock(regs_64_clock),
    .reset(regs_64_reset),
    .io_in(regs_64_io_in),
    .io_init(regs_64_io_init),
    .io_reset(regs_64_io_reset),
    .io_out(regs_64_io_out),
    .io_enable(regs_64_io_enable)
  );
  FF_136 regs_65 (
    .clock(regs_65_clock),
    .reset(regs_65_reset),
    .io_in(regs_65_io_in),
    .io_init(regs_65_io_init),
    .io_reset(regs_65_io_reset),
    .io_out(regs_65_io_out),
    .io_enable(regs_65_io_enable)
  );
  FF_136 regs_66 (
    .clock(regs_66_clock),
    .reset(regs_66_reset),
    .io_in(regs_66_io_in),
    .io_init(regs_66_io_init),
    .io_reset(regs_66_io_reset),
    .io_out(regs_66_io_out),
    .io_enable(regs_66_io_enable)
  );
  FF_136 regs_67 (
    .clock(regs_67_clock),
    .reset(regs_67_reset),
    .io_in(regs_67_io_in),
    .io_init(regs_67_io_init),
    .io_reset(regs_67_io_reset),
    .io_out(regs_67_io_out),
    .io_enable(regs_67_io_enable)
  );
  FF_136 regs_68 (
    .clock(regs_68_clock),
    .reset(regs_68_reset),
    .io_in(regs_68_io_in),
    .io_init(regs_68_io_init),
    .io_reset(regs_68_io_reset),
    .io_out(regs_68_io_out),
    .io_enable(regs_68_io_enable)
  );
  FF_136 regs_69 (
    .clock(regs_69_clock),
    .reset(regs_69_reset),
    .io_in(regs_69_io_in),
    .io_init(regs_69_io_init),
    .io_reset(regs_69_io_reset),
    .io_out(regs_69_io_out),
    .io_enable(regs_69_io_enable)
  );
  FF_136 regs_70 (
    .clock(regs_70_clock),
    .reset(regs_70_reset),
    .io_in(regs_70_io_in),
    .io_init(regs_70_io_init),
    .io_reset(regs_70_io_reset),
    .io_out(regs_70_io_out),
    .io_enable(regs_70_io_enable)
  );
  FF_136 regs_71 (
    .clock(regs_71_clock),
    .reset(regs_71_reset),
    .io_in(regs_71_io_in),
    .io_init(regs_71_io_init),
    .io_reset(regs_71_io_reset),
    .io_out(regs_71_io_out),
    .io_enable(regs_71_io_enable)
  );
  FF_136 regs_72 (
    .clock(regs_72_clock),
    .reset(regs_72_reset),
    .io_in(regs_72_io_in),
    .io_init(regs_72_io_init),
    .io_reset(regs_72_io_reset),
    .io_out(regs_72_io_out),
    .io_enable(regs_72_io_enable)
  );
  FF_136 regs_73 (
    .clock(regs_73_clock),
    .reset(regs_73_reset),
    .io_in(regs_73_io_in),
    .io_init(regs_73_io_init),
    .io_reset(regs_73_io_reset),
    .io_out(regs_73_io_out),
    .io_enable(regs_73_io_enable)
  );
  FF_136 regs_74 (
    .clock(regs_74_clock),
    .reset(regs_74_reset),
    .io_in(regs_74_io_in),
    .io_init(regs_74_io_init),
    .io_reset(regs_74_io_reset),
    .io_out(regs_74_io_out),
    .io_enable(regs_74_io_enable)
  );
  FF_136 regs_75 (
    .clock(regs_75_clock),
    .reset(regs_75_reset),
    .io_in(regs_75_io_in),
    .io_init(regs_75_io_init),
    .io_reset(regs_75_io_reset),
    .io_out(regs_75_io_out),
    .io_enable(regs_75_io_enable)
  );
  FF_136 regs_76 (
    .clock(regs_76_clock),
    .reset(regs_76_reset),
    .io_in(regs_76_io_in),
    .io_init(regs_76_io_init),
    .io_reset(regs_76_io_reset),
    .io_out(regs_76_io_out),
    .io_enable(regs_76_io_enable)
  );
  FF_136 regs_77 (
    .clock(regs_77_clock),
    .reset(regs_77_reset),
    .io_in(regs_77_io_in),
    .io_init(regs_77_io_init),
    .io_reset(regs_77_io_reset),
    .io_out(regs_77_io_out),
    .io_enable(regs_77_io_enable)
  );
  FF_136 regs_78 (
    .clock(regs_78_clock),
    .reset(regs_78_reset),
    .io_in(regs_78_io_in),
    .io_init(regs_78_io_init),
    .io_reset(regs_78_io_reset),
    .io_out(regs_78_io_out),
    .io_enable(regs_78_io_enable)
  );
  FF_136 regs_79 (
    .clock(regs_79_clock),
    .reset(regs_79_reset),
    .io_in(regs_79_io_in),
    .io_init(regs_79_io_init),
    .io_reset(regs_79_io_reset),
    .io_out(regs_79_io_out),
    .io_enable(regs_79_io_enable)
  );
  FF_136 regs_80 (
    .clock(regs_80_clock),
    .reset(regs_80_reset),
    .io_in(regs_80_io_in),
    .io_init(regs_80_io_init),
    .io_reset(regs_80_io_reset),
    .io_out(regs_80_io_out),
    .io_enable(regs_80_io_enable)
  );
  FF_136 regs_81 (
    .clock(regs_81_clock),
    .reset(regs_81_reset),
    .io_in(regs_81_io_in),
    .io_init(regs_81_io_init),
    .io_reset(regs_81_io_reset),
    .io_out(regs_81_io_out),
    .io_enable(regs_81_io_enable)
  );
  FF_136 regs_82 (
    .clock(regs_82_clock),
    .reset(regs_82_reset),
    .io_in(regs_82_io_in),
    .io_init(regs_82_io_init),
    .io_reset(regs_82_io_reset),
    .io_out(regs_82_io_out),
    .io_enable(regs_82_io_enable)
  );
  FF_136 regs_83 (
    .clock(regs_83_clock),
    .reset(regs_83_reset),
    .io_in(regs_83_io_in),
    .io_init(regs_83_io_init),
    .io_reset(regs_83_io_reset),
    .io_out(regs_83_io_out),
    .io_enable(regs_83_io_enable)
  );
  FF_136 regs_84 (
    .clock(regs_84_clock),
    .reset(regs_84_reset),
    .io_in(regs_84_io_in),
    .io_init(regs_84_io_init),
    .io_reset(regs_84_io_reset),
    .io_out(regs_84_io_out),
    .io_enable(regs_84_io_enable)
  );
  FF_136 regs_85 (
    .clock(regs_85_clock),
    .reset(regs_85_reset),
    .io_in(regs_85_io_in),
    .io_init(regs_85_io_init),
    .io_reset(regs_85_io_reset),
    .io_out(regs_85_io_out),
    .io_enable(regs_85_io_enable)
  );
  FF_136 regs_86 (
    .clock(regs_86_clock),
    .reset(regs_86_reset),
    .io_in(regs_86_io_in),
    .io_init(regs_86_io_init),
    .io_reset(regs_86_io_reset),
    .io_out(regs_86_io_out),
    .io_enable(regs_86_io_enable)
  );
  FF_136 regs_87 (
    .clock(regs_87_clock),
    .reset(regs_87_reset),
    .io_in(regs_87_io_in),
    .io_init(regs_87_io_init),
    .io_reset(regs_87_io_reset),
    .io_out(regs_87_io_out),
    .io_enable(regs_87_io_enable)
  );
  FF_136 regs_88 (
    .clock(regs_88_clock),
    .reset(regs_88_reset),
    .io_in(regs_88_io_in),
    .io_init(regs_88_io_init),
    .io_reset(regs_88_io_reset),
    .io_out(regs_88_io_out),
    .io_enable(regs_88_io_enable)
  );
  FF_136 regs_89 (
    .clock(regs_89_clock),
    .reset(regs_89_reset),
    .io_in(regs_89_io_in),
    .io_init(regs_89_io_init),
    .io_reset(regs_89_io_reset),
    .io_out(regs_89_io_out),
    .io_enable(regs_89_io_enable)
  );
  FF_136 regs_90 (
    .clock(regs_90_clock),
    .reset(regs_90_reset),
    .io_in(regs_90_io_in),
    .io_init(regs_90_io_init),
    .io_reset(regs_90_io_reset),
    .io_out(regs_90_io_out),
    .io_enable(regs_90_io_enable)
  );
  FF_136 regs_91 (
    .clock(regs_91_clock),
    .reset(regs_91_reset),
    .io_in(regs_91_io_in),
    .io_init(regs_91_io_init),
    .io_reset(regs_91_io_reset),
    .io_out(regs_91_io_out),
    .io_enable(regs_91_io_enable)
  );
  FF_136 regs_92 (
    .clock(regs_92_clock),
    .reset(regs_92_reset),
    .io_in(regs_92_io_in),
    .io_init(regs_92_io_init),
    .io_reset(regs_92_io_reset),
    .io_out(regs_92_io_out),
    .io_enable(regs_92_io_enable)
  );
  FF_136 regs_93 (
    .clock(regs_93_clock),
    .reset(regs_93_reset),
    .io_in(regs_93_io_in),
    .io_init(regs_93_io_init),
    .io_reset(regs_93_io_reset),
    .io_out(regs_93_io_out),
    .io_enable(regs_93_io_enable)
  );
  FF_136 regs_94 (
    .clock(regs_94_clock),
    .reset(regs_94_reset),
    .io_in(regs_94_io_in),
    .io_init(regs_94_io_init),
    .io_reset(regs_94_io_reset),
    .io_out(regs_94_io_out),
    .io_enable(regs_94_io_enable)
  );
  FF_136 regs_95 (
    .clock(regs_95_clock),
    .reset(regs_95_reset),
    .io_in(regs_95_io_in),
    .io_init(regs_95_io_init),
    .io_reset(regs_95_io_reset),
    .io_out(regs_95_io_out),
    .io_enable(regs_95_io_enable)
  );
  FF_136 regs_96 (
    .clock(regs_96_clock),
    .reset(regs_96_reset),
    .io_in(regs_96_io_in),
    .io_init(regs_96_io_init),
    .io_reset(regs_96_io_reset),
    .io_out(regs_96_io_out),
    .io_enable(regs_96_io_enable)
  );
  FF_136 regs_97 (
    .clock(regs_97_clock),
    .reset(regs_97_reset),
    .io_in(regs_97_io_in),
    .io_init(regs_97_io_init),
    .io_reset(regs_97_io_reset),
    .io_out(regs_97_io_out),
    .io_enable(regs_97_io_enable)
  );
  FF_136 regs_98 (
    .clock(regs_98_clock),
    .reset(regs_98_reset),
    .io_in(regs_98_io_in),
    .io_init(regs_98_io_init),
    .io_reset(regs_98_io_reset),
    .io_out(regs_98_io_out),
    .io_enable(regs_98_io_enable)
  );
  FF_136 regs_99 (
    .clock(regs_99_clock),
    .reset(regs_99_reset),
    .io_in(regs_99_io_in),
    .io_init(regs_99_io_init),
    .io_reset(regs_99_io_reset),
    .io_out(regs_99_io_out),
    .io_enable(regs_99_io_enable)
  );
  FF_136 regs_100 (
    .clock(regs_100_clock),
    .reset(regs_100_reset),
    .io_in(regs_100_io_in),
    .io_init(regs_100_io_init),
    .io_reset(regs_100_io_reset),
    .io_out(regs_100_io_out),
    .io_enable(regs_100_io_enable)
  );
  FF_136 regs_101 (
    .clock(regs_101_clock),
    .reset(regs_101_reset),
    .io_in(regs_101_io_in),
    .io_init(regs_101_io_init),
    .io_reset(regs_101_io_reset),
    .io_out(regs_101_io_out),
    .io_enable(regs_101_io_enable)
  );
  FF_136 regs_102 (
    .clock(regs_102_clock),
    .reset(regs_102_reset),
    .io_in(regs_102_io_in),
    .io_init(regs_102_io_init),
    .io_reset(regs_102_io_reset),
    .io_out(regs_102_io_out),
    .io_enable(regs_102_io_enable)
  );
  FF_136 regs_103 (
    .clock(regs_103_clock),
    .reset(regs_103_reset),
    .io_in(regs_103_io_in),
    .io_init(regs_103_io_init),
    .io_reset(regs_103_io_reset),
    .io_out(regs_103_io_out),
    .io_enable(regs_103_io_enable)
  );
  FF_136 regs_104 (
    .clock(regs_104_clock),
    .reset(regs_104_reset),
    .io_in(regs_104_io_in),
    .io_init(regs_104_io_init),
    .io_reset(regs_104_io_reset),
    .io_out(regs_104_io_out),
    .io_enable(regs_104_io_enable)
  );
  FF_136 regs_105 (
    .clock(regs_105_clock),
    .reset(regs_105_reset),
    .io_in(regs_105_io_in),
    .io_init(regs_105_io_init),
    .io_reset(regs_105_io_reset),
    .io_out(regs_105_io_out),
    .io_enable(regs_105_io_enable)
  );
  FF_136 regs_106 (
    .clock(regs_106_clock),
    .reset(regs_106_reset),
    .io_in(regs_106_io_in),
    .io_init(regs_106_io_init),
    .io_reset(regs_106_io_reset),
    .io_out(regs_106_io_out),
    .io_enable(regs_106_io_enable)
  );
  FF_136 regs_107 (
    .clock(regs_107_clock),
    .reset(regs_107_reset),
    .io_in(regs_107_io_in),
    .io_init(regs_107_io_init),
    .io_reset(regs_107_io_reset),
    .io_out(regs_107_io_out),
    .io_enable(regs_107_io_enable)
  );
  FF_136 regs_108 (
    .clock(regs_108_clock),
    .reset(regs_108_reset),
    .io_in(regs_108_io_in),
    .io_init(regs_108_io_init),
    .io_reset(regs_108_io_reset),
    .io_out(regs_108_io_out),
    .io_enable(regs_108_io_enable)
  );
  FF_136 regs_109 (
    .clock(regs_109_clock),
    .reset(regs_109_reset),
    .io_in(regs_109_io_in),
    .io_init(regs_109_io_init),
    .io_reset(regs_109_io_reset),
    .io_out(regs_109_io_out),
    .io_enable(regs_109_io_enable)
  );
  FF_136 regs_110 (
    .clock(regs_110_clock),
    .reset(regs_110_reset),
    .io_in(regs_110_io_in),
    .io_init(regs_110_io_init),
    .io_reset(regs_110_io_reset),
    .io_out(regs_110_io_out),
    .io_enable(regs_110_io_enable)
  );
  FF_136 regs_111 (
    .clock(regs_111_clock),
    .reset(regs_111_reset),
    .io_in(regs_111_io_in),
    .io_init(regs_111_io_init),
    .io_reset(regs_111_io_reset),
    .io_out(regs_111_io_out),
    .io_enable(regs_111_io_enable)
  );
  FF_136 regs_112 (
    .clock(regs_112_clock),
    .reset(regs_112_reset),
    .io_in(regs_112_io_in),
    .io_init(regs_112_io_init),
    .io_reset(regs_112_io_reset),
    .io_out(regs_112_io_out),
    .io_enable(regs_112_io_enable)
  );
  FF_136 regs_113 (
    .clock(regs_113_clock),
    .reset(regs_113_reset),
    .io_in(regs_113_io_in),
    .io_init(regs_113_io_init),
    .io_reset(regs_113_io_reset),
    .io_out(regs_113_io_out),
    .io_enable(regs_113_io_enable)
  );
  FF_136 regs_114 (
    .clock(regs_114_clock),
    .reset(regs_114_reset),
    .io_in(regs_114_io_in),
    .io_init(regs_114_io_init),
    .io_reset(regs_114_io_reset),
    .io_out(regs_114_io_out),
    .io_enable(regs_114_io_enable)
  );
  FF_136 regs_115 (
    .clock(regs_115_clock),
    .reset(regs_115_reset),
    .io_in(regs_115_io_in),
    .io_init(regs_115_io_init),
    .io_reset(regs_115_io_reset),
    .io_out(regs_115_io_out),
    .io_enable(regs_115_io_enable)
  );
  FF_136 regs_116 (
    .clock(regs_116_clock),
    .reset(regs_116_reset),
    .io_in(regs_116_io_in),
    .io_init(regs_116_io_init),
    .io_reset(regs_116_io_reset),
    .io_out(regs_116_io_out),
    .io_enable(regs_116_io_enable)
  );
  FF_136 regs_117 (
    .clock(regs_117_clock),
    .reset(regs_117_reset),
    .io_in(regs_117_io_in),
    .io_init(regs_117_io_init),
    .io_reset(regs_117_io_reset),
    .io_out(regs_117_io_out),
    .io_enable(regs_117_io_enable)
  );
  FF_136 regs_118 (
    .clock(regs_118_clock),
    .reset(regs_118_reset),
    .io_in(regs_118_io_in),
    .io_init(regs_118_io_init),
    .io_reset(regs_118_io_reset),
    .io_out(regs_118_io_out),
    .io_enable(regs_118_io_enable)
  );
  FF_136 regs_119 (
    .clock(regs_119_clock),
    .reset(regs_119_reset),
    .io_in(regs_119_io_in),
    .io_init(regs_119_io_init),
    .io_reset(regs_119_io_reset),
    .io_out(regs_119_io_out),
    .io_enable(regs_119_io_enable)
  );
  FF_136 regs_120 (
    .clock(regs_120_clock),
    .reset(regs_120_reset),
    .io_in(regs_120_io_in),
    .io_init(regs_120_io_init),
    .io_reset(regs_120_io_reset),
    .io_out(regs_120_io_out),
    .io_enable(regs_120_io_enable)
  );
  FF_136 regs_121 (
    .clock(regs_121_clock),
    .reset(regs_121_reset),
    .io_in(regs_121_io_in),
    .io_init(regs_121_io_init),
    .io_reset(regs_121_io_reset),
    .io_out(regs_121_io_out),
    .io_enable(regs_121_io_enable)
  );
  FF_136 regs_122 (
    .clock(regs_122_clock),
    .reset(regs_122_reset),
    .io_in(regs_122_io_in),
    .io_init(regs_122_io_init),
    .io_reset(regs_122_io_reset),
    .io_out(regs_122_io_out),
    .io_enable(regs_122_io_enable)
  );
  FF_136 regs_123 (
    .clock(regs_123_clock),
    .reset(regs_123_reset),
    .io_in(regs_123_io_in),
    .io_init(regs_123_io_init),
    .io_reset(regs_123_io_reset),
    .io_out(regs_123_io_out),
    .io_enable(regs_123_io_enable)
  );
  FF_136 regs_124 (
    .clock(regs_124_clock),
    .reset(regs_124_reset),
    .io_in(regs_124_io_in),
    .io_init(regs_124_io_init),
    .io_reset(regs_124_io_reset),
    .io_out(regs_124_io_out),
    .io_enable(regs_124_io_enable)
  );
  FF_136 regs_125 (
    .clock(regs_125_clock),
    .reset(regs_125_reset),
    .io_in(regs_125_io_in),
    .io_init(regs_125_io_init),
    .io_reset(regs_125_io_reset),
    .io_out(regs_125_io_out),
    .io_enable(regs_125_io_enable)
  );
  FF_136 regs_126 (
    .clock(regs_126_clock),
    .reset(regs_126_reset),
    .io_in(regs_126_io_in),
    .io_init(regs_126_io_init),
    .io_reset(regs_126_io_reset),
    .io_out(regs_126_io_out),
    .io_enable(regs_126_io_enable)
  );
  FF_136 regs_127 (
    .clock(regs_127_clock),
    .reset(regs_127_reset),
    .io_in(regs_127_io_in),
    .io_init(regs_127_io_init),
    .io_reset(regs_127_io_reset),
    .io_out(regs_127_io_out),
    .io_enable(regs_127_io_enable)
  );
  FF_136 regs_128 (
    .clock(regs_128_clock),
    .reset(regs_128_reset),
    .io_in(regs_128_io_in),
    .io_init(regs_128_io_init),
    .io_reset(regs_128_io_reset),
    .io_out(regs_128_io_out),
    .io_enable(regs_128_io_enable)
  );
  FF_136 regs_129 (
    .clock(regs_129_clock),
    .reset(regs_129_reset),
    .io_in(regs_129_io_in),
    .io_init(regs_129_io_init),
    .io_reset(regs_129_io_reset),
    .io_out(regs_129_io_out),
    .io_enable(regs_129_io_enable)
  );
  FF_136 regs_130 (
    .clock(regs_130_clock),
    .reset(regs_130_reset),
    .io_in(regs_130_io_in),
    .io_init(regs_130_io_init),
    .io_reset(regs_130_io_reset),
    .io_out(regs_130_io_out),
    .io_enable(regs_130_io_enable)
  );
  FF_136 regs_131 (
    .clock(regs_131_clock),
    .reset(regs_131_reset),
    .io_in(regs_131_io_in),
    .io_init(regs_131_io_init),
    .io_reset(regs_131_io_reset),
    .io_out(regs_131_io_out),
    .io_enable(regs_131_io_enable)
  );
  FF_136 regs_132 (
    .clock(regs_132_clock),
    .reset(regs_132_reset),
    .io_in(regs_132_io_in),
    .io_init(regs_132_io_init),
    .io_reset(regs_132_io_reset),
    .io_out(regs_132_io_out),
    .io_enable(regs_132_io_enable)
  );
  FF_136 regs_133 (
    .clock(regs_133_clock),
    .reset(regs_133_reset),
    .io_in(regs_133_io_in),
    .io_init(regs_133_io_init),
    .io_reset(regs_133_io_reset),
    .io_out(regs_133_io_out),
    .io_enable(regs_133_io_enable)
  );
  FF_136 regs_134 (
    .clock(regs_134_clock),
    .reset(regs_134_reset),
    .io_in(regs_134_io_in),
    .io_init(regs_134_io_init),
    .io_reset(regs_134_io_reset),
    .io_out(regs_134_io_out),
    .io_enable(regs_134_io_enable)
  );
  FF_136 regs_135 (
    .clock(regs_135_clock),
    .reset(regs_135_reset),
    .io_in(regs_135_io_in),
    .io_init(regs_135_io_init),
    .io_reset(regs_135_io_reset),
    .io_out(regs_135_io_out),
    .io_enable(regs_135_io_enable)
  );
  FF_136 regs_136 (
    .clock(regs_136_clock),
    .reset(regs_136_reset),
    .io_in(regs_136_io_in),
    .io_init(regs_136_io_init),
    .io_reset(regs_136_io_reset),
    .io_out(regs_136_io_out),
    .io_enable(regs_136_io_enable)
  );
  FF_136 regs_137 (
    .clock(regs_137_clock),
    .reset(regs_137_reset),
    .io_in(regs_137_io_in),
    .io_init(regs_137_io_init),
    .io_reset(regs_137_io_reset),
    .io_out(regs_137_io_out),
    .io_enable(regs_137_io_enable)
  );
  FF_136 regs_138 (
    .clock(regs_138_clock),
    .reset(regs_138_reset),
    .io_in(regs_138_io_in),
    .io_init(regs_138_io_init),
    .io_reset(regs_138_io_reset),
    .io_out(regs_138_io_out),
    .io_enable(regs_138_io_enable)
  );
  FF_136 regs_139 (
    .clock(regs_139_clock),
    .reset(regs_139_reset),
    .io_in(regs_139_io_in),
    .io_init(regs_139_io_init),
    .io_reset(regs_139_io_reset),
    .io_out(regs_139_io_out),
    .io_enable(regs_139_io_enable)
  );
  FF_136 regs_140 (
    .clock(regs_140_clock),
    .reset(regs_140_reset),
    .io_in(regs_140_io_in),
    .io_init(regs_140_io_init),
    .io_reset(regs_140_io_reset),
    .io_out(regs_140_io_out),
    .io_enable(regs_140_io_enable)
  );
  FF_136 regs_141 (
    .clock(regs_141_clock),
    .reset(regs_141_reset),
    .io_in(regs_141_io_in),
    .io_init(regs_141_io_init),
    .io_reset(regs_141_io_reset),
    .io_out(regs_141_io_out),
    .io_enable(regs_141_io_enable)
  );
  FF_136 regs_142 (
    .clock(regs_142_clock),
    .reset(regs_142_reset),
    .io_in(regs_142_io_in),
    .io_init(regs_142_io_init),
    .io_reset(regs_142_io_reset),
    .io_out(regs_142_io_out),
    .io_enable(regs_142_io_enable)
  );
  FF_136 regs_143 (
    .clock(regs_143_clock),
    .reset(regs_143_reset),
    .io_in(regs_143_io_in),
    .io_init(regs_143_io_init),
    .io_reset(regs_143_io_reset),
    .io_out(regs_143_io_out),
    .io_enable(regs_143_io_enable)
  );
  FF_136 regs_144 (
    .clock(regs_144_clock),
    .reset(regs_144_reset),
    .io_in(regs_144_io_in),
    .io_init(regs_144_io_init),
    .io_reset(regs_144_io_reset),
    .io_out(regs_144_io_out),
    .io_enable(regs_144_io_enable)
  );
  FF_136 regs_145 (
    .clock(regs_145_clock),
    .reset(regs_145_reset),
    .io_in(regs_145_io_in),
    .io_init(regs_145_io_init),
    .io_reset(regs_145_io_reset),
    .io_out(regs_145_io_out),
    .io_enable(regs_145_io_enable)
  );
  FF_136 regs_146 (
    .clock(regs_146_clock),
    .reset(regs_146_reset),
    .io_in(regs_146_io_in),
    .io_init(regs_146_io_init),
    .io_reset(regs_146_io_reset),
    .io_out(regs_146_io_out),
    .io_enable(regs_146_io_enable)
  );
  FF_136 regs_147 (
    .clock(regs_147_clock),
    .reset(regs_147_reset),
    .io_in(regs_147_io_in),
    .io_init(regs_147_io_init),
    .io_reset(regs_147_io_reset),
    .io_out(regs_147_io_out),
    .io_enable(regs_147_io_enable)
  );
  FF_136 regs_148 (
    .clock(regs_148_clock),
    .reset(regs_148_reset),
    .io_in(regs_148_io_in),
    .io_init(regs_148_io_init),
    .io_reset(regs_148_io_reset),
    .io_out(regs_148_io_out),
    .io_enable(regs_148_io_enable)
  );
  FF_136 regs_149 (
    .clock(regs_149_clock),
    .reset(regs_149_reset),
    .io_in(regs_149_io_in),
    .io_init(regs_149_io_init),
    .io_reset(regs_149_io_reset),
    .io_out(regs_149_io_out),
    .io_enable(regs_149_io_enable)
  );
  FF_136 regs_150 (
    .clock(regs_150_clock),
    .reset(regs_150_reset),
    .io_in(regs_150_io_in),
    .io_init(regs_150_io_init),
    .io_reset(regs_150_io_reset),
    .io_out(regs_150_io_out),
    .io_enable(regs_150_io_enable)
  );
  FF_136 regs_151 (
    .clock(regs_151_clock),
    .reset(regs_151_reset),
    .io_in(regs_151_io_in),
    .io_init(regs_151_io_init),
    .io_reset(regs_151_io_reset),
    .io_out(regs_151_io_out),
    .io_enable(regs_151_io_enable)
  );
  FF_136 regs_152 (
    .clock(regs_152_clock),
    .reset(regs_152_reset),
    .io_in(regs_152_io_in),
    .io_init(regs_152_io_init),
    .io_reset(regs_152_io_reset),
    .io_out(regs_152_io_out),
    .io_enable(regs_152_io_enable)
  );
  FF_136 regs_153 (
    .clock(regs_153_clock),
    .reset(regs_153_reset),
    .io_in(regs_153_io_in),
    .io_init(regs_153_io_init),
    .io_reset(regs_153_io_reset),
    .io_out(regs_153_io_out),
    .io_enable(regs_153_io_enable)
  );
  FF_136 regs_154 (
    .clock(regs_154_clock),
    .reset(regs_154_reset),
    .io_in(regs_154_io_in),
    .io_init(regs_154_io_init),
    .io_reset(regs_154_io_reset),
    .io_out(regs_154_io_out),
    .io_enable(regs_154_io_enable)
  );
  FF_136 regs_155 (
    .clock(regs_155_clock),
    .reset(regs_155_reset),
    .io_in(regs_155_io_in),
    .io_init(regs_155_io_init),
    .io_reset(regs_155_io_reset),
    .io_out(regs_155_io_out),
    .io_enable(regs_155_io_enable)
  );
  FF_136 regs_156 (
    .clock(regs_156_clock),
    .reset(regs_156_reset),
    .io_in(regs_156_io_in),
    .io_init(regs_156_io_init),
    .io_reset(regs_156_io_reset),
    .io_out(regs_156_io_out),
    .io_enable(regs_156_io_enable)
  );
  FF_136 regs_157 (
    .clock(regs_157_clock),
    .reset(regs_157_reset),
    .io_in(regs_157_io_in),
    .io_init(regs_157_io_init),
    .io_reset(regs_157_io_reset),
    .io_out(regs_157_io_out),
    .io_enable(regs_157_io_enable)
  );
  FF_136 regs_158 (
    .clock(regs_158_clock),
    .reset(regs_158_reset),
    .io_in(regs_158_io_in),
    .io_init(regs_158_io_init),
    .io_reset(regs_158_io_reset),
    .io_out(regs_158_io_out),
    .io_enable(regs_158_io_enable)
  );
  FF_136 regs_159 (
    .clock(regs_159_clock),
    .reset(regs_159_reset),
    .io_in(regs_159_io_in),
    .io_init(regs_159_io_init),
    .io_reset(regs_159_io_reset),
    .io_out(regs_159_io_out),
    .io_enable(regs_159_io_enable)
  );
  FF_136 regs_160 (
    .clock(regs_160_clock),
    .reset(regs_160_reset),
    .io_in(regs_160_io_in),
    .io_init(regs_160_io_init),
    .io_reset(regs_160_io_reset),
    .io_out(regs_160_io_out),
    .io_enable(regs_160_io_enable)
  );
  FF_136 regs_161 (
    .clock(regs_161_clock),
    .reset(regs_161_reset),
    .io_in(regs_161_io_in),
    .io_init(regs_161_io_init),
    .io_reset(regs_161_io_reset),
    .io_out(regs_161_io_out),
    .io_enable(regs_161_io_enable)
  );
  FF_136 regs_162 (
    .clock(regs_162_clock),
    .reset(regs_162_reset),
    .io_in(regs_162_io_in),
    .io_init(regs_162_io_init),
    .io_reset(regs_162_io_reset),
    .io_out(regs_162_io_out),
    .io_enable(regs_162_io_enable)
  );
  FF_136 regs_163 (
    .clock(regs_163_clock),
    .reset(regs_163_reset),
    .io_in(regs_163_io_in),
    .io_init(regs_163_io_init),
    .io_reset(regs_163_io_reset),
    .io_out(regs_163_io_out),
    .io_enable(regs_163_io_enable)
  );
  FF_136 regs_164 (
    .clock(regs_164_clock),
    .reset(regs_164_reset),
    .io_in(regs_164_io_in),
    .io_init(regs_164_io_init),
    .io_reset(regs_164_io_reset),
    .io_out(regs_164_io_out),
    .io_enable(regs_164_io_enable)
  );
  FF_136 regs_165 (
    .clock(regs_165_clock),
    .reset(regs_165_reset),
    .io_in(regs_165_io_in),
    .io_init(regs_165_io_init),
    .io_reset(regs_165_io_reset),
    .io_out(regs_165_io_out),
    .io_enable(regs_165_io_enable)
  );
  FF_136 regs_166 (
    .clock(regs_166_clock),
    .reset(regs_166_reset),
    .io_in(regs_166_io_in),
    .io_init(regs_166_io_init),
    .io_reset(regs_166_io_reset),
    .io_out(regs_166_io_out),
    .io_enable(regs_166_io_enable)
  );
  FF_136 regs_167 (
    .clock(regs_167_clock),
    .reset(regs_167_reset),
    .io_in(regs_167_io_in),
    .io_init(regs_167_io_init),
    .io_reset(regs_167_io_reset),
    .io_out(regs_167_io_out),
    .io_enable(regs_167_io_enable)
  );
  FF_136 regs_168 (
    .clock(regs_168_clock),
    .reset(regs_168_reset),
    .io_in(regs_168_io_in),
    .io_init(regs_168_io_init),
    .io_reset(regs_168_io_reset),
    .io_out(regs_168_io_out),
    .io_enable(regs_168_io_enable)
  );
  FF_136 regs_169 (
    .clock(regs_169_clock),
    .reset(regs_169_reset),
    .io_in(regs_169_io_in),
    .io_init(regs_169_io_init),
    .io_reset(regs_169_io_reset),
    .io_out(regs_169_io_out),
    .io_enable(regs_169_io_enable)
  );
  FF_136 regs_170 (
    .clock(regs_170_clock),
    .reset(regs_170_reset),
    .io_in(regs_170_io_in),
    .io_init(regs_170_io_init),
    .io_reset(regs_170_io_reset),
    .io_out(regs_170_io_out),
    .io_enable(regs_170_io_enable)
  );
  FF_136 regs_171 (
    .clock(regs_171_clock),
    .reset(regs_171_reset),
    .io_in(regs_171_io_in),
    .io_init(regs_171_io_init),
    .io_reset(regs_171_io_reset),
    .io_out(regs_171_io_out),
    .io_enable(regs_171_io_enable)
  );
  FF_136 regs_172 (
    .clock(regs_172_clock),
    .reset(regs_172_reset),
    .io_in(regs_172_io_in),
    .io_init(regs_172_io_init),
    .io_reset(regs_172_io_reset),
    .io_out(regs_172_io_out),
    .io_enable(regs_172_io_enable)
  );
  FF_136 regs_173 (
    .clock(regs_173_clock),
    .reset(regs_173_reset),
    .io_in(regs_173_io_in),
    .io_init(regs_173_io_init),
    .io_reset(regs_173_io_reset),
    .io_out(regs_173_io_out),
    .io_enable(regs_173_io_enable)
  );
  FF_136 regs_174 (
    .clock(regs_174_clock),
    .reset(regs_174_reset),
    .io_in(regs_174_io_in),
    .io_init(regs_174_io_init),
    .io_reset(regs_174_io_reset),
    .io_out(regs_174_io_out),
    .io_enable(regs_174_io_enable)
  );
  FF_136 regs_175 (
    .clock(regs_175_clock),
    .reset(regs_175_reset),
    .io_in(regs_175_io_in),
    .io_init(regs_175_io_init),
    .io_reset(regs_175_io_reset),
    .io_out(regs_175_io_out),
    .io_enable(regs_175_io_enable)
  );
  FF_136 regs_176 (
    .clock(regs_176_clock),
    .reset(regs_176_reset),
    .io_in(regs_176_io_in),
    .io_init(regs_176_io_init),
    .io_reset(regs_176_io_reset),
    .io_out(regs_176_io_out),
    .io_enable(regs_176_io_enable)
  );
  FF_136 regs_177 (
    .clock(regs_177_clock),
    .reset(regs_177_reset),
    .io_in(regs_177_io_in),
    .io_init(regs_177_io_init),
    .io_reset(regs_177_io_reset),
    .io_out(regs_177_io_out),
    .io_enable(regs_177_io_enable)
  );
  FF_136 regs_178 (
    .clock(regs_178_clock),
    .reset(regs_178_reset),
    .io_in(regs_178_io_in),
    .io_init(regs_178_io_init),
    .io_reset(regs_178_io_reset),
    .io_out(regs_178_io_out),
    .io_enable(regs_178_io_enable)
  );
  FF_136 regs_179 (
    .clock(regs_179_clock),
    .reset(regs_179_reset),
    .io_in(regs_179_io_in),
    .io_init(regs_179_io_init),
    .io_reset(regs_179_io_reset),
    .io_out(regs_179_io_out),
    .io_enable(regs_179_io_enable)
  );
  FF_136 regs_180 (
    .clock(regs_180_clock),
    .reset(regs_180_reset),
    .io_in(regs_180_io_in),
    .io_init(regs_180_io_init),
    .io_reset(regs_180_io_reset),
    .io_out(regs_180_io_out),
    .io_enable(regs_180_io_enable)
  );
  FF_136 regs_181 (
    .clock(regs_181_clock),
    .reset(regs_181_reset),
    .io_in(regs_181_io_in),
    .io_init(regs_181_io_init),
    .io_reset(regs_181_io_reset),
    .io_out(regs_181_io_out),
    .io_enable(regs_181_io_enable)
  );
  FF_136 regs_182 (
    .clock(regs_182_clock),
    .reset(regs_182_reset),
    .io_in(regs_182_io_in),
    .io_init(regs_182_io_init),
    .io_reset(regs_182_io_reset),
    .io_out(regs_182_io_out),
    .io_enable(regs_182_io_enable)
  );
  FF_136 regs_183 (
    .clock(regs_183_clock),
    .reset(regs_183_reset),
    .io_in(regs_183_io_in),
    .io_init(regs_183_io_init),
    .io_reset(regs_183_io_reset),
    .io_out(regs_183_io_out),
    .io_enable(regs_183_io_enable)
  );
  FF_136 regs_184 (
    .clock(regs_184_clock),
    .reset(regs_184_reset),
    .io_in(regs_184_io_in),
    .io_init(regs_184_io_init),
    .io_reset(regs_184_io_reset),
    .io_out(regs_184_io_out),
    .io_enable(regs_184_io_enable)
  );
  FF_136 regs_185 (
    .clock(regs_185_clock),
    .reset(regs_185_reset),
    .io_in(regs_185_io_in),
    .io_init(regs_185_io_init),
    .io_reset(regs_185_io_reset),
    .io_out(regs_185_io_out),
    .io_enable(regs_185_io_enable)
  );
  FF_136 regs_186 (
    .clock(regs_186_clock),
    .reset(regs_186_reset),
    .io_in(regs_186_io_in),
    .io_init(regs_186_io_init),
    .io_reset(regs_186_io_reset),
    .io_out(regs_186_io_out),
    .io_enable(regs_186_io_enable)
  );
  FF_136 regs_187 (
    .clock(regs_187_clock),
    .reset(regs_187_reset),
    .io_in(regs_187_io_in),
    .io_init(regs_187_io_init),
    .io_reset(regs_187_io_reset),
    .io_out(regs_187_io_out),
    .io_enable(regs_187_io_enable)
  );
  FF_136 regs_188 (
    .clock(regs_188_clock),
    .reset(regs_188_reset),
    .io_in(regs_188_io_in),
    .io_init(regs_188_io_init),
    .io_reset(regs_188_io_reset),
    .io_out(regs_188_io_out),
    .io_enable(regs_188_io_enable)
  );
  FF_136 regs_189 (
    .clock(regs_189_clock),
    .reset(regs_189_reset),
    .io_in(regs_189_io_in),
    .io_init(regs_189_io_init),
    .io_reset(regs_189_io_reset),
    .io_out(regs_189_io_out),
    .io_enable(regs_189_io_enable)
  );
  FF_136 regs_190 (
    .clock(regs_190_clock),
    .reset(regs_190_reset),
    .io_in(regs_190_io_in),
    .io_init(regs_190_io_init),
    .io_reset(regs_190_io_reset),
    .io_out(regs_190_io_out),
    .io_enable(regs_190_io_enable)
  );
  FF_136 regs_191 (
    .clock(regs_191_clock),
    .reset(regs_191_reset),
    .io_in(regs_191_io_in),
    .io_init(regs_191_io_init),
    .io_reset(regs_191_io_reset),
    .io_out(regs_191_io_out),
    .io_enable(regs_191_io_enable)
  );
  FF_136 regs_192 (
    .clock(regs_192_clock),
    .reset(regs_192_reset),
    .io_in(regs_192_io_in),
    .io_init(regs_192_io_init),
    .io_reset(regs_192_io_reset),
    .io_out(regs_192_io_out),
    .io_enable(regs_192_io_enable)
  );
  FF_136 regs_193 (
    .clock(regs_193_clock),
    .reset(regs_193_reset),
    .io_in(regs_193_io_in),
    .io_init(regs_193_io_init),
    .io_reset(regs_193_io_reset),
    .io_out(regs_193_io_out),
    .io_enable(regs_193_io_enable)
  );
  FF_136 regs_194 (
    .clock(regs_194_clock),
    .reset(regs_194_reset),
    .io_in(regs_194_io_in),
    .io_init(regs_194_io_init),
    .io_reset(regs_194_io_reset),
    .io_out(regs_194_io_out),
    .io_enable(regs_194_io_enable)
  );
  FF_136 regs_195 (
    .clock(regs_195_clock),
    .reset(regs_195_reset),
    .io_in(regs_195_io_in),
    .io_init(regs_195_io_init),
    .io_reset(regs_195_io_reset),
    .io_out(regs_195_io_out),
    .io_enable(regs_195_io_enable)
  );
  FF_136 regs_196 (
    .clock(regs_196_clock),
    .reset(regs_196_reset),
    .io_in(regs_196_io_in),
    .io_init(regs_196_io_init),
    .io_reset(regs_196_io_reset),
    .io_out(regs_196_io_out),
    .io_enable(regs_196_io_enable)
  );
  FF_136 regs_197 (
    .clock(regs_197_clock),
    .reset(regs_197_reset),
    .io_in(regs_197_io_in),
    .io_init(regs_197_io_init),
    .io_reset(regs_197_io_reset),
    .io_out(regs_197_io_out),
    .io_enable(regs_197_io_enable)
  );
  FF_136 regs_198 (
    .clock(regs_198_clock),
    .reset(regs_198_reset),
    .io_in(regs_198_io_in),
    .io_init(regs_198_io_init),
    .io_reset(regs_198_io_reset),
    .io_out(regs_198_io_out),
    .io_enable(regs_198_io_enable)
  );
  FF_136 regs_199 (
    .clock(regs_199_clock),
    .reset(regs_199_reset),
    .io_in(regs_199_io_in),
    .io_init(regs_199_io_init),
    .io_reset(regs_199_io_reset),
    .io_out(regs_199_io_out),
    .io_enable(regs_199_io_enable)
  );
  FF_136 regs_200 (
    .clock(regs_200_clock),
    .reset(regs_200_reset),
    .io_in(regs_200_io_in),
    .io_init(regs_200_io_init),
    .io_reset(regs_200_io_reset),
    .io_out(regs_200_io_out),
    .io_enable(regs_200_io_enable)
  );
  FF_136 regs_201 (
    .clock(regs_201_clock),
    .reset(regs_201_reset),
    .io_in(regs_201_io_in),
    .io_init(regs_201_io_init),
    .io_reset(regs_201_io_reset),
    .io_out(regs_201_io_out),
    .io_enable(regs_201_io_enable)
  );
  FF_136 regs_202 (
    .clock(regs_202_clock),
    .reset(regs_202_reset),
    .io_in(regs_202_io_in),
    .io_init(regs_202_io_init),
    .io_reset(regs_202_io_reset),
    .io_out(regs_202_io_out),
    .io_enable(regs_202_io_enable)
  );
  FF_136 regs_203 (
    .clock(regs_203_clock),
    .reset(regs_203_reset),
    .io_in(regs_203_io_in),
    .io_init(regs_203_io_init),
    .io_reset(regs_203_io_reset),
    .io_out(regs_203_io_out),
    .io_enable(regs_203_io_enable)
  );
  FF_136 regs_204 (
    .clock(regs_204_clock),
    .reset(regs_204_reset),
    .io_in(regs_204_io_in),
    .io_init(regs_204_io_init),
    .io_reset(regs_204_io_reset),
    .io_out(regs_204_io_out),
    .io_enable(regs_204_io_enable)
  );
  FF_136 regs_205 (
    .clock(regs_205_clock),
    .reset(regs_205_reset),
    .io_in(regs_205_io_in),
    .io_init(regs_205_io_init),
    .io_reset(regs_205_io_reset),
    .io_out(regs_205_io_out),
    .io_enable(regs_205_io_enable)
  );
  FF_136 regs_206 (
    .clock(regs_206_clock),
    .reset(regs_206_reset),
    .io_in(regs_206_io_in),
    .io_init(regs_206_io_init),
    .io_reset(regs_206_io_reset),
    .io_out(regs_206_io_out),
    .io_enable(regs_206_io_enable)
  );
  FF_136 regs_207 (
    .clock(regs_207_clock),
    .reset(regs_207_reset),
    .io_in(regs_207_io_in),
    .io_init(regs_207_io_init),
    .io_reset(regs_207_io_reset),
    .io_out(regs_207_io_out),
    .io_enable(regs_207_io_enable)
  );
  FF_136 regs_208 (
    .clock(regs_208_clock),
    .reset(regs_208_reset),
    .io_in(regs_208_io_in),
    .io_init(regs_208_io_init),
    .io_reset(regs_208_io_reset),
    .io_out(regs_208_io_out),
    .io_enable(regs_208_io_enable)
  );
  FF_136 regs_209 (
    .clock(regs_209_clock),
    .reset(regs_209_reset),
    .io_in(regs_209_io_in),
    .io_init(regs_209_io_init),
    .io_reset(regs_209_io_reset),
    .io_out(regs_209_io_out),
    .io_enable(regs_209_io_enable)
  );
  FF_136 regs_210 (
    .clock(regs_210_clock),
    .reset(regs_210_reset),
    .io_in(regs_210_io_in),
    .io_init(regs_210_io_init),
    .io_reset(regs_210_io_reset),
    .io_out(regs_210_io_out),
    .io_enable(regs_210_io_enable)
  );
  FF_136 regs_211 (
    .clock(regs_211_clock),
    .reset(regs_211_reset),
    .io_in(regs_211_io_in),
    .io_init(regs_211_io_init),
    .io_reset(regs_211_io_reset),
    .io_out(regs_211_io_out),
    .io_enable(regs_211_io_enable)
  );
  FF_136 regs_212 (
    .clock(regs_212_clock),
    .reset(regs_212_reset),
    .io_in(regs_212_io_in),
    .io_init(regs_212_io_init),
    .io_reset(regs_212_io_reset),
    .io_out(regs_212_io_out),
    .io_enable(regs_212_io_enable)
  );
  FF_136 regs_213 (
    .clock(regs_213_clock),
    .reset(regs_213_reset),
    .io_in(regs_213_io_in),
    .io_init(regs_213_io_init),
    .io_reset(regs_213_io_reset),
    .io_out(regs_213_io_out),
    .io_enable(regs_213_io_enable)
  );
  FF_136 regs_214 (
    .clock(regs_214_clock),
    .reset(regs_214_reset),
    .io_in(regs_214_io_in),
    .io_init(regs_214_io_init),
    .io_reset(regs_214_io_reset),
    .io_out(regs_214_io_out),
    .io_enable(regs_214_io_enable)
  );
  FF_136 regs_215 (
    .clock(regs_215_clock),
    .reset(regs_215_reset),
    .io_in(regs_215_io_in),
    .io_init(regs_215_io_init),
    .io_reset(regs_215_io_reset),
    .io_out(regs_215_io_out),
    .io_enable(regs_215_io_enable)
  );
  FF_136 regs_216 (
    .clock(regs_216_clock),
    .reset(regs_216_reset),
    .io_in(regs_216_io_in),
    .io_init(regs_216_io_init),
    .io_reset(regs_216_io_reset),
    .io_out(regs_216_io_out),
    .io_enable(regs_216_io_enable)
  );
  FF_136 regs_217 (
    .clock(regs_217_clock),
    .reset(regs_217_reset),
    .io_in(regs_217_io_in),
    .io_init(regs_217_io_init),
    .io_reset(regs_217_io_reset),
    .io_out(regs_217_io_out),
    .io_enable(regs_217_io_enable)
  );
  FF_136 regs_218 (
    .clock(regs_218_clock),
    .reset(regs_218_reset),
    .io_in(regs_218_io_in),
    .io_init(regs_218_io_init),
    .io_reset(regs_218_io_reset),
    .io_out(regs_218_io_out),
    .io_enable(regs_218_io_enable)
  );
  FF_136 regs_219 (
    .clock(regs_219_clock),
    .reset(regs_219_reset),
    .io_in(regs_219_io_in),
    .io_init(regs_219_io_init),
    .io_reset(regs_219_io_reset),
    .io_out(regs_219_io_out),
    .io_enable(regs_219_io_enable)
  );
  FF_136 regs_220 (
    .clock(regs_220_clock),
    .reset(regs_220_reset),
    .io_in(regs_220_io_in),
    .io_init(regs_220_io_init),
    .io_reset(regs_220_io_reset),
    .io_out(regs_220_io_out),
    .io_enable(regs_220_io_enable)
  );
  FF_136 regs_221 (
    .clock(regs_221_clock),
    .reset(regs_221_reset),
    .io_in(regs_221_io_in),
    .io_init(regs_221_io_init),
    .io_reset(regs_221_io_reset),
    .io_out(regs_221_io_out),
    .io_enable(regs_221_io_enable)
  );
  FF_136 regs_222 (
    .clock(regs_222_clock),
    .reset(regs_222_reset),
    .io_in(regs_222_io_in),
    .io_init(regs_222_io_init),
    .io_reset(regs_222_io_reset),
    .io_out(regs_222_io_out),
    .io_enable(regs_222_io_enable)
  );
  FF_136 regs_223 (
    .clock(regs_223_clock),
    .reset(regs_223_reset),
    .io_in(regs_223_io_in),
    .io_init(regs_223_io_init),
    .io_reset(regs_223_io_reset),
    .io_out(regs_223_io_out),
    .io_enable(regs_223_io_enable)
  );
  FF_136 regs_224 (
    .clock(regs_224_clock),
    .reset(regs_224_reset),
    .io_in(regs_224_io_in),
    .io_init(regs_224_io_init),
    .io_reset(regs_224_io_reset),
    .io_out(regs_224_io_out),
    .io_enable(regs_224_io_enable)
  );
  FF_136 regs_225 (
    .clock(regs_225_clock),
    .reset(regs_225_reset),
    .io_in(regs_225_io_in),
    .io_init(regs_225_io_init),
    .io_reset(regs_225_io_reset),
    .io_out(regs_225_io_out),
    .io_enable(regs_225_io_enable)
  );
  FF_136 regs_226 (
    .clock(regs_226_clock),
    .reset(regs_226_reset),
    .io_in(regs_226_io_in),
    .io_init(regs_226_io_init),
    .io_reset(regs_226_io_reset),
    .io_out(regs_226_io_out),
    .io_enable(regs_226_io_enable)
  );
  FF_136 regs_227 (
    .clock(regs_227_clock),
    .reset(regs_227_reset),
    .io_in(regs_227_io_in),
    .io_init(regs_227_io_init),
    .io_reset(regs_227_io_reset),
    .io_out(regs_227_io_out),
    .io_enable(regs_227_io_enable)
  );
  FF_136 regs_228 (
    .clock(regs_228_clock),
    .reset(regs_228_reset),
    .io_in(regs_228_io_in),
    .io_init(regs_228_io_init),
    .io_reset(regs_228_io_reset),
    .io_out(regs_228_io_out),
    .io_enable(regs_228_io_enable)
  );
  FF_136 regs_229 (
    .clock(regs_229_clock),
    .reset(regs_229_reset),
    .io_in(regs_229_io_in),
    .io_init(regs_229_io_init),
    .io_reset(regs_229_io_reset),
    .io_out(regs_229_io_out),
    .io_enable(regs_229_io_enable)
  );
  FF_136 regs_230 (
    .clock(regs_230_clock),
    .reset(regs_230_reset),
    .io_in(regs_230_io_in),
    .io_init(regs_230_io_init),
    .io_reset(regs_230_io_reset),
    .io_out(regs_230_io_out),
    .io_enable(regs_230_io_enable)
  );
  FF_136 regs_231 (
    .clock(regs_231_clock),
    .reset(regs_231_reset),
    .io_in(regs_231_io_in),
    .io_init(regs_231_io_init),
    .io_reset(regs_231_io_reset),
    .io_out(regs_231_io_out),
    .io_enable(regs_231_io_enable)
  );
  FF_136 regs_232 (
    .clock(regs_232_clock),
    .reset(regs_232_reset),
    .io_in(regs_232_io_in),
    .io_init(regs_232_io_init),
    .io_reset(regs_232_io_reset),
    .io_out(regs_232_io_out),
    .io_enable(regs_232_io_enable)
  );
  FF_136 regs_233 (
    .clock(regs_233_clock),
    .reset(regs_233_reset),
    .io_in(regs_233_io_in),
    .io_init(regs_233_io_init),
    .io_reset(regs_233_io_reset),
    .io_out(regs_233_io_out),
    .io_enable(regs_233_io_enable)
  );
  FF_136 regs_234 (
    .clock(regs_234_clock),
    .reset(regs_234_reset),
    .io_in(regs_234_io_in),
    .io_init(regs_234_io_init),
    .io_reset(regs_234_io_reset),
    .io_out(regs_234_io_out),
    .io_enable(regs_234_io_enable)
  );
  FF_136 regs_235 (
    .clock(regs_235_clock),
    .reset(regs_235_reset),
    .io_in(regs_235_io_in),
    .io_init(regs_235_io_init),
    .io_reset(regs_235_io_reset),
    .io_out(regs_235_io_out),
    .io_enable(regs_235_io_enable)
  );
  FF_136 regs_236 (
    .clock(regs_236_clock),
    .reset(regs_236_reset),
    .io_in(regs_236_io_in),
    .io_init(regs_236_io_init),
    .io_reset(regs_236_io_reset),
    .io_out(regs_236_io_out),
    .io_enable(regs_236_io_enable)
  );
  FF_136 regs_237 (
    .clock(regs_237_clock),
    .reset(regs_237_reset),
    .io_in(regs_237_io_in),
    .io_init(regs_237_io_init),
    .io_reset(regs_237_io_reset),
    .io_out(regs_237_io_out),
    .io_enable(regs_237_io_enable)
  );
  FF_136 regs_238 (
    .clock(regs_238_clock),
    .reset(regs_238_reset),
    .io_in(regs_238_io_in),
    .io_init(regs_238_io_init),
    .io_reset(regs_238_io_reset),
    .io_out(regs_238_io_out),
    .io_enable(regs_238_io_enable)
  );
  FF_136 regs_239 (
    .clock(regs_239_clock),
    .reset(regs_239_reset),
    .io_in(regs_239_io_in),
    .io_init(regs_239_io_init),
    .io_reset(regs_239_io_reset),
    .io_out(regs_239_io_out),
    .io_enable(regs_239_io_enable)
  );
  FF_136 regs_240 (
    .clock(regs_240_clock),
    .reset(regs_240_reset),
    .io_in(regs_240_io_in),
    .io_init(regs_240_io_init),
    .io_reset(regs_240_io_reset),
    .io_out(regs_240_io_out),
    .io_enable(regs_240_io_enable)
  );
  FF_136 regs_241 (
    .clock(regs_241_clock),
    .reset(regs_241_reset),
    .io_in(regs_241_io_in),
    .io_init(regs_241_io_init),
    .io_reset(regs_241_io_reset),
    .io_out(regs_241_io_out),
    .io_enable(regs_241_io_enable)
  );
  FF_136 regs_242 (
    .clock(regs_242_clock),
    .reset(regs_242_reset),
    .io_in(regs_242_io_in),
    .io_init(regs_242_io_init),
    .io_reset(regs_242_io_reset),
    .io_out(regs_242_io_out),
    .io_enable(regs_242_io_enable)
  );
  FF_136 regs_243 (
    .clock(regs_243_clock),
    .reset(regs_243_reset),
    .io_in(regs_243_io_in),
    .io_init(regs_243_io_init),
    .io_reset(regs_243_io_reset),
    .io_out(regs_243_io_out),
    .io_enable(regs_243_io_enable)
  );
  FF_136 regs_244 (
    .clock(regs_244_clock),
    .reset(regs_244_reset),
    .io_in(regs_244_io_in),
    .io_init(regs_244_io_init),
    .io_reset(regs_244_io_reset),
    .io_out(regs_244_io_out),
    .io_enable(regs_244_io_enable)
  );
  FF_136 regs_245 (
    .clock(regs_245_clock),
    .reset(regs_245_reset),
    .io_in(regs_245_io_in),
    .io_init(regs_245_io_init),
    .io_reset(regs_245_io_reset),
    .io_out(regs_245_io_out),
    .io_enable(regs_245_io_enable)
  );
  FF_136 regs_246 (
    .clock(regs_246_clock),
    .reset(regs_246_reset),
    .io_in(regs_246_io_in),
    .io_init(regs_246_io_init),
    .io_reset(regs_246_io_reset),
    .io_out(regs_246_io_out),
    .io_enable(regs_246_io_enable)
  );
  FF_136 regs_247 (
    .clock(regs_247_clock),
    .reset(regs_247_reset),
    .io_in(regs_247_io_in),
    .io_init(regs_247_io_init),
    .io_reset(regs_247_io_reset),
    .io_out(regs_247_io_out),
    .io_enable(regs_247_io_enable)
  );
  FF_136 regs_248 (
    .clock(regs_248_clock),
    .reset(regs_248_reset),
    .io_in(regs_248_io_in),
    .io_init(regs_248_io_init),
    .io_reset(regs_248_io_reset),
    .io_out(regs_248_io_out),
    .io_enable(regs_248_io_enable)
  );
  FF_136 regs_249 (
    .clock(regs_249_clock),
    .reset(regs_249_reset),
    .io_in(regs_249_io_in),
    .io_init(regs_249_io_init),
    .io_reset(regs_249_io_reset),
    .io_out(regs_249_io_out),
    .io_enable(regs_249_io_enable)
  );
  FF_136 regs_250 (
    .clock(regs_250_clock),
    .reset(regs_250_reset),
    .io_in(regs_250_io_in),
    .io_init(regs_250_io_init),
    .io_reset(regs_250_io_reset),
    .io_out(regs_250_io_out),
    .io_enable(regs_250_io_enable)
  );
  FF_136 regs_251 (
    .clock(regs_251_clock),
    .reset(regs_251_reset),
    .io_in(regs_251_io_in),
    .io_init(regs_251_io_init),
    .io_reset(regs_251_io_reset),
    .io_out(regs_251_io_out),
    .io_enable(regs_251_io_enable)
  );
  FF_136 regs_252 (
    .clock(regs_252_clock),
    .reset(regs_252_reset),
    .io_in(regs_252_io_in),
    .io_init(regs_252_io_init),
    .io_reset(regs_252_io_reset),
    .io_out(regs_252_io_out),
    .io_enable(regs_252_io_enable)
  );
  FF_136 regs_253 (
    .clock(regs_253_clock),
    .reset(regs_253_reset),
    .io_in(regs_253_io_in),
    .io_init(regs_253_io_init),
    .io_reset(regs_253_io_reset),
    .io_out(regs_253_io_out),
    .io_enable(regs_253_io_enable)
  );
  FF_136 regs_254 (
    .clock(regs_254_clock),
    .reset(regs_254_reset),
    .io_in(regs_254_io_in),
    .io_init(regs_254_io_init),
    .io_reset(regs_254_io_reset),
    .io_out(regs_254_io_out),
    .io_enable(regs_254_io_enable)
  );
  FF_136 regs_255 (
    .clock(regs_255_clock),
    .reset(regs_255_reset),
    .io_in(regs_255_io_in),
    .io_init(regs_255_io_init),
    .io_reset(regs_255_io_reset),
    .io_out(regs_255_io_out),
    .io_enable(regs_255_io_enable)
  );
  FF_136 regs_256 (
    .clock(regs_256_clock),
    .reset(regs_256_reset),
    .io_in(regs_256_io_in),
    .io_init(regs_256_io_init),
    .io_reset(regs_256_io_reset),
    .io_out(regs_256_io_out),
    .io_enable(regs_256_io_enable)
  );
  FF_136 regs_257 (
    .clock(regs_257_clock),
    .reset(regs_257_reset),
    .io_in(regs_257_io_in),
    .io_init(regs_257_io_init),
    .io_reset(regs_257_io_reset),
    .io_out(regs_257_io_out),
    .io_enable(regs_257_io_enable)
  );
  FF_136 regs_258 (
    .clock(regs_258_clock),
    .reset(regs_258_reset),
    .io_in(regs_258_io_in),
    .io_init(regs_258_io_init),
    .io_reset(regs_258_io_reset),
    .io_out(regs_258_io_out),
    .io_enable(regs_258_io_enable)
  );
  FF_136 regs_259 (
    .clock(regs_259_clock),
    .reset(regs_259_reset),
    .io_in(regs_259_io_in),
    .io_init(regs_259_io_init),
    .io_reset(regs_259_io_reset),
    .io_out(regs_259_io_out),
    .io_enable(regs_259_io_enable)
  );
  FF_136 regs_260 (
    .clock(regs_260_clock),
    .reset(regs_260_reset),
    .io_in(regs_260_io_in),
    .io_init(regs_260_io_init),
    .io_reset(regs_260_io_reset),
    .io_out(regs_260_io_out),
    .io_enable(regs_260_io_enable)
  );
  FF_136 regs_261 (
    .clock(regs_261_clock),
    .reset(regs_261_reset),
    .io_in(regs_261_io_in),
    .io_init(regs_261_io_init),
    .io_reset(regs_261_io_reset),
    .io_out(regs_261_io_out),
    .io_enable(regs_261_io_enable)
  );
  FF_136 regs_262 (
    .clock(regs_262_clock),
    .reset(regs_262_reset),
    .io_in(regs_262_io_in),
    .io_init(regs_262_io_init),
    .io_reset(regs_262_io_reset),
    .io_out(regs_262_io_out),
    .io_enable(regs_262_io_enable)
  );
  FF_136 regs_263 (
    .clock(regs_263_clock),
    .reset(regs_263_reset),
    .io_in(regs_263_io_in),
    .io_init(regs_263_io_init),
    .io_reset(regs_263_io_reset),
    .io_out(regs_263_io_out),
    .io_enable(regs_263_io_enable)
  );
  FF_136 regs_264 (
    .clock(regs_264_clock),
    .reset(regs_264_reset),
    .io_in(regs_264_io_in),
    .io_init(regs_264_io_init),
    .io_reset(regs_264_io_reset),
    .io_out(regs_264_io_out),
    .io_enable(regs_264_io_enable)
  );
  FF_136 regs_265 (
    .clock(regs_265_clock),
    .reset(regs_265_reset),
    .io_in(regs_265_io_in),
    .io_init(regs_265_io_init),
    .io_reset(regs_265_io_reset),
    .io_out(regs_265_io_out),
    .io_enable(regs_265_io_enable)
  );
  FF_136 regs_266 (
    .clock(regs_266_clock),
    .reset(regs_266_reset),
    .io_in(regs_266_io_in),
    .io_init(regs_266_io_init),
    .io_reset(regs_266_io_reset),
    .io_out(regs_266_io_out),
    .io_enable(regs_266_io_enable)
  );
  FF_136 regs_267 (
    .clock(regs_267_clock),
    .reset(regs_267_reset),
    .io_in(regs_267_io_in),
    .io_init(regs_267_io_init),
    .io_reset(regs_267_io_reset),
    .io_out(regs_267_io_out),
    .io_enable(regs_267_io_enable)
  );
  FF_136 regs_268 (
    .clock(regs_268_clock),
    .reset(regs_268_reset),
    .io_in(regs_268_io_in),
    .io_init(regs_268_io_init),
    .io_reset(regs_268_io_reset),
    .io_out(regs_268_io_out),
    .io_enable(regs_268_io_enable)
  );
  FF_136 regs_269 (
    .clock(regs_269_clock),
    .reset(regs_269_reset),
    .io_in(regs_269_io_in),
    .io_init(regs_269_io_init),
    .io_reset(regs_269_io_reset),
    .io_out(regs_269_io_out),
    .io_enable(regs_269_io_enable)
  );
  FF_136 regs_270 (
    .clock(regs_270_clock),
    .reset(regs_270_reset),
    .io_in(regs_270_io_in),
    .io_init(regs_270_io_init),
    .io_reset(regs_270_io_reset),
    .io_out(regs_270_io_out),
    .io_enable(regs_270_io_enable)
  );
  FF_136 regs_271 (
    .clock(regs_271_clock),
    .reset(regs_271_reset),
    .io_in(regs_271_io_in),
    .io_init(regs_271_io_init),
    .io_reset(regs_271_io_reset),
    .io_out(regs_271_io_out),
    .io_enable(regs_271_io_enable)
  );
  FF_136 regs_272 (
    .clock(regs_272_clock),
    .reset(regs_272_reset),
    .io_in(regs_272_io_in),
    .io_init(regs_272_io_init),
    .io_reset(regs_272_io_reset),
    .io_out(regs_272_io_out),
    .io_enable(regs_272_io_enable)
  );
  FF_136 regs_273 (
    .clock(regs_273_clock),
    .reset(regs_273_reset),
    .io_in(regs_273_io_in),
    .io_init(regs_273_io_init),
    .io_reset(regs_273_io_reset),
    .io_out(regs_273_io_out),
    .io_enable(regs_273_io_enable)
  );
  FF_136 regs_274 (
    .clock(regs_274_clock),
    .reset(regs_274_reset),
    .io_in(regs_274_io_in),
    .io_init(regs_274_io_init),
    .io_reset(regs_274_io_reset),
    .io_out(regs_274_io_out),
    .io_enable(regs_274_io_enable)
  );
  FF_136 regs_275 (
    .clock(regs_275_clock),
    .reset(regs_275_reset),
    .io_in(regs_275_io_in),
    .io_init(regs_275_io_init),
    .io_reset(regs_275_io_reset),
    .io_out(regs_275_io_out),
    .io_enable(regs_275_io_enable)
  );
  FF_136 regs_276 (
    .clock(regs_276_clock),
    .reset(regs_276_reset),
    .io_in(regs_276_io_in),
    .io_init(regs_276_io_init),
    .io_reset(regs_276_io_reset),
    .io_out(regs_276_io_out),
    .io_enable(regs_276_io_enable)
  );
  FF_136 regs_277 (
    .clock(regs_277_clock),
    .reset(regs_277_reset),
    .io_in(regs_277_io_in),
    .io_init(regs_277_io_init),
    .io_reset(regs_277_io_reset),
    .io_out(regs_277_io_out),
    .io_enable(regs_277_io_enable)
  );
  FF_136 regs_278 (
    .clock(regs_278_clock),
    .reset(regs_278_reset),
    .io_in(regs_278_io_in),
    .io_init(regs_278_io_init),
    .io_reset(regs_278_io_reset),
    .io_out(regs_278_io_out),
    .io_enable(regs_278_io_enable)
  );
  FF_136 regs_279 (
    .clock(regs_279_clock),
    .reset(regs_279_reset),
    .io_in(regs_279_io_in),
    .io_init(regs_279_io_init),
    .io_reset(regs_279_io_reset),
    .io_out(regs_279_io_out),
    .io_enable(regs_279_io_enable)
  );
  FF_136 regs_280 (
    .clock(regs_280_clock),
    .reset(regs_280_reset),
    .io_in(regs_280_io_in),
    .io_init(regs_280_io_init),
    .io_reset(regs_280_io_reset),
    .io_out(regs_280_io_out),
    .io_enable(regs_280_io_enable)
  );
  FF_136 regs_281 (
    .clock(regs_281_clock),
    .reset(regs_281_reset),
    .io_in(regs_281_io_in),
    .io_init(regs_281_io_init),
    .io_reset(regs_281_io_reset),
    .io_out(regs_281_io_out),
    .io_enable(regs_281_io_enable)
  );
  FF_136 regs_282 (
    .clock(regs_282_clock),
    .reset(regs_282_reset),
    .io_in(regs_282_io_in),
    .io_init(regs_282_io_init),
    .io_reset(regs_282_io_reset),
    .io_out(regs_282_io_out),
    .io_enable(regs_282_io_enable)
  );
  FF_136 regs_283 (
    .clock(regs_283_clock),
    .reset(regs_283_reset),
    .io_in(regs_283_io_in),
    .io_init(regs_283_io_init),
    .io_reset(regs_283_io_reset),
    .io_out(regs_283_io_out),
    .io_enable(regs_283_io_enable)
  );
  FF_136 regs_284 (
    .clock(regs_284_clock),
    .reset(regs_284_reset),
    .io_in(regs_284_io_in),
    .io_init(regs_284_io_init),
    .io_reset(regs_284_io_reset),
    .io_out(regs_284_io_out),
    .io_enable(regs_284_io_enable)
  );
  FF_136 regs_285 (
    .clock(regs_285_clock),
    .reset(regs_285_reset),
    .io_in(regs_285_io_in),
    .io_init(regs_285_io_init),
    .io_reset(regs_285_io_reset),
    .io_out(regs_285_io_out),
    .io_enable(regs_285_io_enable)
  );
  FF_136 regs_286 (
    .clock(regs_286_clock),
    .reset(regs_286_reset),
    .io_in(regs_286_io_in),
    .io_init(regs_286_io_init),
    .io_reset(regs_286_io_reset),
    .io_out(regs_286_io_out),
    .io_enable(regs_286_io_enable)
  );
  FF_136 regs_287 (
    .clock(regs_287_clock),
    .reset(regs_287_reset),
    .io_in(regs_287_io_in),
    .io_init(regs_287_io_init),
    .io_reset(regs_287_io_reset),
    .io_out(regs_287_io_out),
    .io_enable(regs_287_io_enable)
  );
  FF_136 regs_288 (
    .clock(regs_288_clock),
    .reset(regs_288_reset),
    .io_in(regs_288_io_in),
    .io_init(regs_288_io_init),
    .io_reset(regs_288_io_reset),
    .io_out(regs_288_io_out),
    .io_enable(regs_288_io_enable)
  );
  FF_136 regs_289 (
    .clock(regs_289_clock),
    .reset(regs_289_reset),
    .io_in(regs_289_io_in),
    .io_init(regs_289_io_init),
    .io_reset(regs_289_io_reset),
    .io_out(regs_289_io_out),
    .io_enable(regs_289_io_enable)
  );
  FF_136 regs_290 (
    .clock(regs_290_clock),
    .reset(regs_290_reset),
    .io_in(regs_290_io_in),
    .io_init(regs_290_io_init),
    .io_reset(regs_290_io_reset),
    .io_out(regs_290_io_out),
    .io_enable(regs_290_io_enable)
  );
  FF_136 regs_291 (
    .clock(regs_291_clock),
    .reset(regs_291_reset),
    .io_in(regs_291_io_in),
    .io_init(regs_291_io_init),
    .io_reset(regs_291_io_reset),
    .io_out(regs_291_io_out),
    .io_enable(regs_291_io_enable)
  );
  FF_136 regs_292 (
    .clock(regs_292_clock),
    .reset(regs_292_reset),
    .io_in(regs_292_io_in),
    .io_init(regs_292_io_init),
    .io_reset(regs_292_io_reset),
    .io_out(regs_292_io_out),
    .io_enable(regs_292_io_enable)
  );
  FF_136 regs_293 (
    .clock(regs_293_clock),
    .reset(regs_293_reset),
    .io_in(regs_293_io_in),
    .io_init(regs_293_io_init),
    .io_reset(regs_293_io_reset),
    .io_out(regs_293_io_out),
    .io_enable(regs_293_io_enable)
  );
  FF_136 regs_294 (
    .clock(regs_294_clock),
    .reset(regs_294_reset),
    .io_in(regs_294_io_in),
    .io_init(regs_294_io_init),
    .io_reset(regs_294_io_reset),
    .io_out(regs_294_io_out),
    .io_enable(regs_294_io_enable)
  );
  FF_136 regs_295 (
    .clock(regs_295_clock),
    .reset(regs_295_reset),
    .io_in(regs_295_io_in),
    .io_init(regs_295_io_init),
    .io_reset(regs_295_io_reset),
    .io_out(regs_295_io_out),
    .io_enable(regs_295_io_enable)
  );
  FF_136 regs_296 (
    .clock(regs_296_clock),
    .reset(regs_296_reset),
    .io_in(regs_296_io_in),
    .io_init(regs_296_io_init),
    .io_reset(regs_296_io_reset),
    .io_out(regs_296_io_out),
    .io_enable(regs_296_io_enable)
  );
  FF_136 regs_297 (
    .clock(regs_297_clock),
    .reset(regs_297_reset),
    .io_in(regs_297_io_in),
    .io_init(regs_297_io_init),
    .io_reset(regs_297_io_reset),
    .io_out(regs_297_io_out),
    .io_enable(regs_297_io_enable)
  );
  FF_136 regs_298 (
    .clock(regs_298_clock),
    .reset(regs_298_reset),
    .io_in(regs_298_io_in),
    .io_init(regs_298_io_init),
    .io_reset(regs_298_io_reset),
    .io_out(regs_298_io_out),
    .io_enable(regs_298_io_enable)
  );
  FF_136 regs_299 (
    .clock(regs_299_clock),
    .reset(regs_299_reset),
    .io_in(regs_299_io_in),
    .io_init(regs_299_io_init),
    .io_reset(regs_299_io_reset),
    .io_out(regs_299_io_out),
    .io_enable(regs_299_io_enable)
  );
  FF_136 regs_300 (
    .clock(regs_300_clock),
    .reset(regs_300_reset),
    .io_in(regs_300_io_in),
    .io_init(regs_300_io_init),
    .io_reset(regs_300_io_reset),
    .io_out(regs_300_io_out),
    .io_enable(regs_300_io_enable)
  );
  FF_136 regs_301 (
    .clock(regs_301_clock),
    .reset(regs_301_reset),
    .io_in(regs_301_io_in),
    .io_init(regs_301_io_init),
    .io_reset(regs_301_io_reset),
    .io_out(regs_301_io_out),
    .io_enable(regs_301_io_enable)
  );
  FF_136 regs_302 (
    .clock(regs_302_clock),
    .reset(regs_302_reset),
    .io_in(regs_302_io_in),
    .io_init(regs_302_io_init),
    .io_reset(regs_302_io_reset),
    .io_out(regs_302_io_out),
    .io_enable(regs_302_io_enable)
  );
  FF_136 regs_303 (
    .clock(regs_303_clock),
    .reset(regs_303_reset),
    .io_in(regs_303_io_in),
    .io_init(regs_303_io_init),
    .io_reset(regs_303_io_reset),
    .io_out(regs_303_io_out),
    .io_enable(regs_303_io_enable)
  );
  FF_136 regs_304 (
    .clock(regs_304_clock),
    .reset(regs_304_reset),
    .io_in(regs_304_io_in),
    .io_init(regs_304_io_init),
    .io_reset(regs_304_io_reset),
    .io_out(regs_304_io_out),
    .io_enable(regs_304_io_enable)
  );
  FF_136 regs_305 (
    .clock(regs_305_clock),
    .reset(regs_305_reset),
    .io_in(regs_305_io_in),
    .io_init(regs_305_io_init),
    .io_reset(regs_305_io_reset),
    .io_out(regs_305_io_out),
    .io_enable(regs_305_io_enable)
  );
  FF_136 regs_306 (
    .clock(regs_306_clock),
    .reset(regs_306_reset),
    .io_in(regs_306_io_in),
    .io_init(regs_306_io_init),
    .io_reset(regs_306_io_reset),
    .io_out(regs_306_io_out),
    .io_enable(regs_306_io_enable)
  );
  FF_136 regs_307 (
    .clock(regs_307_clock),
    .reset(regs_307_reset),
    .io_in(regs_307_io_in),
    .io_init(regs_307_io_init),
    .io_reset(regs_307_io_reset),
    .io_out(regs_307_io_out),
    .io_enable(regs_307_io_enable)
  );
  FF_136 regs_308 (
    .clock(regs_308_clock),
    .reset(regs_308_reset),
    .io_in(regs_308_io_in),
    .io_init(regs_308_io_init),
    .io_reset(regs_308_io_reset),
    .io_out(regs_308_io_out),
    .io_enable(regs_308_io_enable)
  );
  FF_136 regs_309 (
    .clock(regs_309_clock),
    .reset(regs_309_reset),
    .io_in(regs_309_io_in),
    .io_init(regs_309_io_init),
    .io_reset(regs_309_io_reset),
    .io_out(regs_309_io_out),
    .io_enable(regs_309_io_enable)
  );
  FF_136 regs_310 (
    .clock(regs_310_clock),
    .reset(regs_310_reset),
    .io_in(regs_310_io_in),
    .io_init(regs_310_io_init),
    .io_reset(regs_310_io_reset),
    .io_out(regs_310_io_out),
    .io_enable(regs_310_io_enable)
  );
  FF_136 regs_311 (
    .clock(regs_311_clock),
    .reset(regs_311_reset),
    .io_in(regs_311_io_in),
    .io_init(regs_311_io_init),
    .io_reset(regs_311_io_reset),
    .io_out(regs_311_io_out),
    .io_enable(regs_311_io_enable)
  );
  FF_136 regs_312 (
    .clock(regs_312_clock),
    .reset(regs_312_reset),
    .io_in(regs_312_io_in),
    .io_init(regs_312_io_init),
    .io_reset(regs_312_io_reset),
    .io_out(regs_312_io_out),
    .io_enable(regs_312_io_enable)
  );
  FF_136 regs_313 (
    .clock(regs_313_clock),
    .reset(regs_313_reset),
    .io_in(regs_313_io_in),
    .io_init(regs_313_io_init),
    .io_reset(regs_313_io_reset),
    .io_out(regs_313_io_out),
    .io_enable(regs_313_io_enable)
  );
  FF_136 regs_314 (
    .clock(regs_314_clock),
    .reset(regs_314_reset),
    .io_in(regs_314_io_in),
    .io_init(regs_314_io_init),
    .io_reset(regs_314_io_reset),
    .io_out(regs_314_io_out),
    .io_enable(regs_314_io_enable)
  );
  FF_136 regs_315 (
    .clock(regs_315_clock),
    .reset(regs_315_reset),
    .io_in(regs_315_io_in),
    .io_init(regs_315_io_init),
    .io_reset(regs_315_io_reset),
    .io_out(regs_315_io_out),
    .io_enable(regs_315_io_enable)
  );
  FF_136 regs_316 (
    .clock(regs_316_clock),
    .reset(regs_316_reset),
    .io_in(regs_316_io_in),
    .io_init(regs_316_io_init),
    .io_reset(regs_316_io_reset),
    .io_out(regs_316_io_out),
    .io_enable(regs_316_io_enable)
  );
  FF_136 regs_317 (
    .clock(regs_317_clock),
    .reset(regs_317_reset),
    .io_in(regs_317_io_in),
    .io_init(regs_317_io_init),
    .io_reset(regs_317_io_reset),
    .io_out(regs_317_io_out),
    .io_enable(regs_317_io_enable)
  );
  FF_136 regs_318 (
    .clock(regs_318_clock),
    .reset(regs_318_reset),
    .io_in(regs_318_io_in),
    .io_init(regs_318_io_init),
    .io_reset(regs_318_io_reset),
    .io_out(regs_318_io_out),
    .io_enable(regs_318_io_enable)
  );
  FF_136 regs_319 (
    .clock(regs_319_clock),
    .reset(regs_319_reset),
    .io_in(regs_319_io_in),
    .io_init(regs_319_io_init),
    .io_reset(regs_319_io_reset),
    .io_out(regs_319_io_out),
    .io_enable(regs_319_io_enable)
  );
  FF_136 regs_320 (
    .clock(regs_320_clock),
    .reset(regs_320_reset),
    .io_in(regs_320_io_in),
    .io_init(regs_320_io_init),
    .io_reset(regs_320_io_reset),
    .io_out(regs_320_io_out),
    .io_enable(regs_320_io_enable)
  );
  FF_136 regs_321 (
    .clock(regs_321_clock),
    .reset(regs_321_reset),
    .io_in(regs_321_io_in),
    .io_init(regs_321_io_init),
    .io_reset(regs_321_io_reset),
    .io_out(regs_321_io_out),
    .io_enable(regs_321_io_enable)
  );
  FF_136 regs_322 (
    .clock(regs_322_clock),
    .reset(regs_322_reset),
    .io_in(regs_322_io_in),
    .io_init(regs_322_io_init),
    .io_reset(regs_322_io_reset),
    .io_out(regs_322_io_out),
    .io_enable(regs_322_io_enable)
  );
  FF_136 regs_323 (
    .clock(regs_323_clock),
    .reset(regs_323_reset),
    .io_in(regs_323_io_in),
    .io_init(regs_323_io_init),
    .io_reset(regs_323_io_reset),
    .io_out(regs_323_io_out),
    .io_enable(regs_323_io_enable)
  );
  FF_136 regs_324 (
    .clock(regs_324_clock),
    .reset(regs_324_reset),
    .io_in(regs_324_io_in),
    .io_init(regs_324_io_init),
    .io_reset(regs_324_io_reset),
    .io_out(regs_324_io_out),
    .io_enable(regs_324_io_enable)
  );
  FF_136 regs_325 (
    .clock(regs_325_clock),
    .reset(regs_325_reset),
    .io_in(regs_325_io_in),
    .io_init(regs_325_io_init),
    .io_reset(regs_325_io_reset),
    .io_out(regs_325_io_out),
    .io_enable(regs_325_io_enable)
  );
  FF_136 regs_326 (
    .clock(regs_326_clock),
    .reset(regs_326_reset),
    .io_in(regs_326_io_in),
    .io_init(regs_326_io_init),
    .io_reset(regs_326_io_reset),
    .io_out(regs_326_io_out),
    .io_enable(regs_326_io_enable)
  );
  FF_136 regs_327 (
    .clock(regs_327_clock),
    .reset(regs_327_reset),
    .io_in(regs_327_io_in),
    .io_init(regs_327_io_init),
    .io_reset(regs_327_io_reset),
    .io_out(regs_327_io_out),
    .io_enable(regs_327_io_enable)
  );
  FF_136 regs_328 (
    .clock(regs_328_clock),
    .reset(regs_328_reset),
    .io_in(regs_328_io_in),
    .io_init(regs_328_io_init),
    .io_reset(regs_328_io_reset),
    .io_out(regs_328_io_out),
    .io_enable(regs_328_io_enable)
  );
  FF_136 regs_329 (
    .clock(regs_329_clock),
    .reset(regs_329_reset),
    .io_in(regs_329_io_in),
    .io_init(regs_329_io_init),
    .io_reset(regs_329_io_reset),
    .io_out(regs_329_io_out),
    .io_enable(regs_329_io_enable)
  );
  FF_136 regs_330 (
    .clock(regs_330_clock),
    .reset(regs_330_reset),
    .io_in(regs_330_io_in),
    .io_init(regs_330_io_init),
    .io_reset(regs_330_io_reset),
    .io_out(regs_330_io_out),
    .io_enable(regs_330_io_enable)
  );
  FF_136 regs_331 (
    .clock(regs_331_clock),
    .reset(regs_331_reset),
    .io_in(regs_331_io_in),
    .io_init(regs_331_io_init),
    .io_reset(regs_331_io_reset),
    .io_out(regs_331_io_out),
    .io_enable(regs_331_io_enable)
  );
  FF_136 regs_332 (
    .clock(regs_332_clock),
    .reset(regs_332_reset),
    .io_in(regs_332_io_in),
    .io_init(regs_332_io_init),
    .io_reset(regs_332_io_reset),
    .io_out(regs_332_io_out),
    .io_enable(regs_332_io_enable)
  );
  FF_136 regs_333 (
    .clock(regs_333_clock),
    .reset(regs_333_reset),
    .io_in(regs_333_io_in),
    .io_init(regs_333_io_init),
    .io_reset(regs_333_io_reset),
    .io_out(regs_333_io_out),
    .io_enable(regs_333_io_enable)
  );
  FF_136 regs_334 (
    .clock(regs_334_clock),
    .reset(regs_334_reset),
    .io_in(regs_334_io_in),
    .io_init(regs_334_io_init),
    .io_reset(regs_334_io_reset),
    .io_out(regs_334_io_out),
    .io_enable(regs_334_io_enable)
  );
  FF_136 regs_335 (
    .clock(regs_335_clock),
    .reset(regs_335_reset),
    .io_in(regs_335_io_in),
    .io_init(regs_335_io_init),
    .io_reset(regs_335_io_reset),
    .io_out(regs_335_io_out),
    .io_enable(regs_335_io_enable)
  );
  FF_136 regs_336 (
    .clock(regs_336_clock),
    .reset(regs_336_reset),
    .io_in(regs_336_io_in),
    .io_init(regs_336_io_init),
    .io_reset(regs_336_io_reset),
    .io_out(regs_336_io_out),
    .io_enable(regs_336_io_enable)
  );
  FF_136 regs_337 (
    .clock(regs_337_clock),
    .reset(regs_337_reset),
    .io_in(regs_337_io_in),
    .io_init(regs_337_io_init),
    .io_reset(regs_337_io_reset),
    .io_out(regs_337_io_out),
    .io_enable(regs_337_io_enable)
  );
  FF_136 regs_338 (
    .clock(regs_338_clock),
    .reset(regs_338_reset),
    .io_in(regs_338_io_in),
    .io_init(regs_338_io_init),
    .io_reset(regs_338_io_reset),
    .io_out(regs_338_io_out),
    .io_enable(regs_338_io_enable)
  );
  FF_136 regs_339 (
    .clock(regs_339_clock),
    .reset(regs_339_reset),
    .io_in(regs_339_io_in),
    .io_init(regs_339_io_init),
    .io_reset(regs_339_io_reset),
    .io_out(regs_339_io_out),
    .io_enable(regs_339_io_enable)
  );
  FF_136 regs_340 (
    .clock(regs_340_clock),
    .reset(regs_340_reset),
    .io_in(regs_340_io_in),
    .io_init(regs_340_io_init),
    .io_reset(regs_340_io_reset),
    .io_out(regs_340_io_out),
    .io_enable(regs_340_io_enable)
  );
  FF_136 regs_341 (
    .clock(regs_341_clock),
    .reset(regs_341_reset),
    .io_in(regs_341_io_in),
    .io_init(regs_341_io_init),
    .io_reset(regs_341_io_reset),
    .io_out(regs_341_io_out),
    .io_enable(regs_341_io_enable)
  );
  FF_136 regs_342 (
    .clock(regs_342_clock),
    .reset(regs_342_reset),
    .io_in(regs_342_io_in),
    .io_init(regs_342_io_init),
    .io_reset(regs_342_io_reset),
    .io_out(regs_342_io_out),
    .io_enable(regs_342_io_enable)
  );
  FF_136 regs_343 (
    .clock(regs_343_clock),
    .reset(regs_343_reset),
    .io_in(regs_343_io_in),
    .io_init(regs_343_io_init),
    .io_reset(regs_343_io_reset),
    .io_out(regs_343_io_out),
    .io_enable(regs_343_io_enable)
  );
  FF_136 regs_344 (
    .clock(regs_344_clock),
    .reset(regs_344_reset),
    .io_in(regs_344_io_in),
    .io_init(regs_344_io_init),
    .io_reset(regs_344_io_reset),
    .io_out(regs_344_io_out),
    .io_enable(regs_344_io_enable)
  );
  FF_136 regs_345 (
    .clock(regs_345_clock),
    .reset(regs_345_reset),
    .io_in(regs_345_io_in),
    .io_init(regs_345_io_init),
    .io_reset(regs_345_io_reset),
    .io_out(regs_345_io_out),
    .io_enable(regs_345_io_enable)
  );
  FF_136 regs_346 (
    .clock(regs_346_clock),
    .reset(regs_346_reset),
    .io_in(regs_346_io_in),
    .io_init(regs_346_io_init),
    .io_reset(regs_346_io_reset),
    .io_out(regs_346_io_out),
    .io_enable(regs_346_io_enable)
  );
  FF_136 regs_347 (
    .clock(regs_347_clock),
    .reset(regs_347_reset),
    .io_in(regs_347_io_in),
    .io_init(regs_347_io_init),
    .io_reset(regs_347_io_reset),
    .io_out(regs_347_io_out),
    .io_enable(regs_347_io_enable)
  );
  FF_136 regs_348 (
    .clock(regs_348_clock),
    .reset(regs_348_reset),
    .io_in(regs_348_io_in),
    .io_init(regs_348_io_init),
    .io_reset(regs_348_io_reset),
    .io_out(regs_348_io_out),
    .io_enable(regs_348_io_enable)
  );
  FF_136 regs_349 (
    .clock(regs_349_clock),
    .reset(regs_349_reset),
    .io_in(regs_349_io_in),
    .io_init(regs_349_io_init),
    .io_reset(regs_349_io_reset),
    .io_out(regs_349_io_out),
    .io_enable(regs_349_io_enable)
  );
  FF_136 regs_350 (
    .clock(regs_350_clock),
    .reset(regs_350_reset),
    .io_in(regs_350_io_in),
    .io_init(regs_350_io_init),
    .io_reset(regs_350_io_reset),
    .io_out(regs_350_io_out),
    .io_enable(regs_350_io_enable)
  );
  FF_136 regs_351 (
    .clock(regs_351_clock),
    .reset(regs_351_reset),
    .io_in(regs_351_io_in),
    .io_init(regs_351_io_init),
    .io_reset(regs_351_io_reset),
    .io_out(regs_351_io_out),
    .io_enable(regs_351_io_enable)
  );
  FF_136 regs_352 (
    .clock(regs_352_clock),
    .reset(regs_352_reset),
    .io_in(regs_352_io_in),
    .io_init(regs_352_io_init),
    .io_reset(regs_352_io_reset),
    .io_out(regs_352_io_out),
    .io_enable(regs_352_io_enable)
  );
  FF_136 regs_353 (
    .clock(regs_353_clock),
    .reset(regs_353_reset),
    .io_in(regs_353_io_in),
    .io_init(regs_353_io_init),
    .io_reset(regs_353_io_reset),
    .io_out(regs_353_io_out),
    .io_enable(regs_353_io_enable)
  );
  FF_136 regs_354 (
    .clock(regs_354_clock),
    .reset(regs_354_reset),
    .io_in(regs_354_io_in),
    .io_init(regs_354_io_init),
    .io_reset(regs_354_io_reset),
    .io_out(regs_354_io_out),
    .io_enable(regs_354_io_enable)
  );
  FF_136 regs_355 (
    .clock(regs_355_clock),
    .reset(regs_355_reset),
    .io_in(regs_355_io_in),
    .io_init(regs_355_io_init),
    .io_reset(regs_355_io_reset),
    .io_out(regs_355_io_out),
    .io_enable(regs_355_io_enable)
  );
  FF_136 regs_356 (
    .clock(regs_356_clock),
    .reset(regs_356_reset),
    .io_in(regs_356_io_in),
    .io_init(regs_356_io_init),
    .io_reset(regs_356_io_reset),
    .io_out(regs_356_io_out),
    .io_enable(regs_356_io_enable)
  );
  FF_136 regs_357 (
    .clock(regs_357_clock),
    .reset(regs_357_reset),
    .io_in(regs_357_io_in),
    .io_init(regs_357_io_init),
    .io_reset(regs_357_io_reset),
    .io_out(regs_357_io_out),
    .io_enable(regs_357_io_enable)
  );
  FF_136 regs_358 (
    .clock(regs_358_clock),
    .reset(regs_358_reset),
    .io_in(regs_358_io_in),
    .io_init(regs_358_io_init),
    .io_reset(regs_358_io_reset),
    .io_out(regs_358_io_out),
    .io_enable(regs_358_io_enable)
  );
  FF_136 regs_359 (
    .clock(regs_359_clock),
    .reset(regs_359_reset),
    .io_in(regs_359_io_in),
    .io_init(regs_359_io_init),
    .io_reset(regs_359_io_reset),
    .io_out(regs_359_io_out),
    .io_enable(regs_359_io_enable)
  );
  FF_136 regs_360 (
    .clock(regs_360_clock),
    .reset(regs_360_reset),
    .io_in(regs_360_io_in),
    .io_init(regs_360_io_init),
    .io_reset(regs_360_io_reset),
    .io_out(regs_360_io_out),
    .io_enable(regs_360_io_enable)
  );
  FF_136 regs_361 (
    .clock(regs_361_clock),
    .reset(regs_361_reset),
    .io_in(regs_361_io_in),
    .io_init(regs_361_io_init),
    .io_reset(regs_361_io_reset),
    .io_out(regs_361_io_out),
    .io_enable(regs_361_io_enable)
  );
  FF_136 regs_362 (
    .clock(regs_362_clock),
    .reset(regs_362_reset),
    .io_in(regs_362_io_in),
    .io_init(regs_362_io_init),
    .io_reset(regs_362_io_reset),
    .io_out(regs_362_io_out),
    .io_enable(regs_362_io_enable)
  );
  FF_136 regs_363 (
    .clock(regs_363_clock),
    .reset(regs_363_reset),
    .io_in(regs_363_io_in),
    .io_init(regs_363_io_init),
    .io_reset(regs_363_io_reset),
    .io_out(regs_363_io_out),
    .io_enable(regs_363_io_enable)
  );
  FF_136 regs_364 (
    .clock(regs_364_clock),
    .reset(regs_364_reset),
    .io_in(regs_364_io_in),
    .io_init(regs_364_io_init),
    .io_reset(regs_364_io_reset),
    .io_out(regs_364_io_out),
    .io_enable(regs_364_io_enable)
  );
  FF_136 regs_365 (
    .clock(regs_365_clock),
    .reset(regs_365_reset),
    .io_in(regs_365_io_in),
    .io_init(regs_365_io_init),
    .io_reset(regs_365_io_reset),
    .io_out(regs_365_io_out),
    .io_enable(regs_365_io_enable)
  );
  FF_136 regs_366 (
    .clock(regs_366_clock),
    .reset(regs_366_reset),
    .io_in(regs_366_io_in),
    .io_init(regs_366_io_init),
    .io_reset(regs_366_io_reset),
    .io_out(regs_366_io_out),
    .io_enable(regs_366_io_enable)
  );
  FF_136 regs_367 (
    .clock(regs_367_clock),
    .reset(regs_367_reset),
    .io_in(regs_367_io_in),
    .io_init(regs_367_io_init),
    .io_reset(regs_367_io_reset),
    .io_out(regs_367_io_out),
    .io_enable(regs_367_io_enable)
  );
  FF_136 regs_368 (
    .clock(regs_368_clock),
    .reset(regs_368_reset),
    .io_in(regs_368_io_in),
    .io_init(regs_368_io_init),
    .io_reset(regs_368_io_reset),
    .io_out(regs_368_io_out),
    .io_enable(regs_368_io_enable)
  );
  FF_136 regs_369 (
    .clock(regs_369_clock),
    .reset(regs_369_reset),
    .io_in(regs_369_io_in),
    .io_init(regs_369_io_init),
    .io_reset(regs_369_io_reset),
    .io_out(regs_369_io_out),
    .io_enable(regs_369_io_enable)
  );
  FF_136 regs_370 (
    .clock(regs_370_clock),
    .reset(regs_370_reset),
    .io_in(regs_370_io_in),
    .io_init(regs_370_io_init),
    .io_reset(regs_370_io_reset),
    .io_out(regs_370_io_out),
    .io_enable(regs_370_io_enable)
  );
  FF_136 regs_371 (
    .clock(regs_371_clock),
    .reset(regs_371_reset),
    .io_in(regs_371_io_in),
    .io_init(regs_371_io_init),
    .io_reset(regs_371_io_reset),
    .io_out(regs_371_io_out),
    .io_enable(regs_371_io_enable)
  );
  FF_136 regs_372 (
    .clock(regs_372_clock),
    .reset(regs_372_reset),
    .io_in(regs_372_io_in),
    .io_init(regs_372_io_init),
    .io_reset(regs_372_io_reset),
    .io_out(regs_372_io_out),
    .io_enable(regs_372_io_enable)
  );
  FF_136 regs_373 (
    .clock(regs_373_clock),
    .reset(regs_373_reset),
    .io_in(regs_373_io_in),
    .io_init(regs_373_io_init),
    .io_reset(regs_373_io_reset),
    .io_out(regs_373_io_out),
    .io_enable(regs_373_io_enable)
  );
  FF_136 regs_374 (
    .clock(regs_374_clock),
    .reset(regs_374_reset),
    .io_in(regs_374_io_in),
    .io_init(regs_374_io_init),
    .io_reset(regs_374_io_reset),
    .io_out(regs_374_io_out),
    .io_enable(regs_374_io_enable)
  );
  FF_136 regs_375 (
    .clock(regs_375_clock),
    .reset(regs_375_reset),
    .io_in(regs_375_io_in),
    .io_init(regs_375_io_init),
    .io_reset(regs_375_io_reset),
    .io_out(regs_375_io_out),
    .io_enable(regs_375_io_enable)
  );
  FF_136 regs_376 (
    .clock(regs_376_clock),
    .reset(regs_376_reset),
    .io_in(regs_376_io_in),
    .io_init(regs_376_io_init),
    .io_reset(regs_376_io_reset),
    .io_out(regs_376_io_out),
    .io_enable(regs_376_io_enable)
  );
  FF_136 regs_377 (
    .clock(regs_377_clock),
    .reset(regs_377_reset),
    .io_in(regs_377_io_in),
    .io_init(regs_377_io_init),
    .io_reset(regs_377_io_reset),
    .io_out(regs_377_io_out),
    .io_enable(regs_377_io_enable)
  );
  FF_136 regs_378 (
    .clock(regs_378_clock),
    .reset(regs_378_reset),
    .io_in(regs_378_io_in),
    .io_init(regs_378_io_init),
    .io_reset(regs_378_io_reset),
    .io_out(regs_378_io_out),
    .io_enable(regs_378_io_enable)
  );
  FF_136 regs_379 (
    .clock(regs_379_clock),
    .reset(regs_379_reset),
    .io_in(regs_379_io_in),
    .io_init(regs_379_io_init),
    .io_reset(regs_379_io_reset),
    .io_out(regs_379_io_out),
    .io_enable(regs_379_io_enable)
  );
  FF_136 regs_380 (
    .clock(regs_380_clock),
    .reset(regs_380_reset),
    .io_in(regs_380_io_in),
    .io_init(regs_380_io_init),
    .io_reset(regs_380_io_reset),
    .io_out(regs_380_io_out),
    .io_enable(regs_380_io_enable)
  );
  FF_136 regs_381 (
    .clock(regs_381_clock),
    .reset(regs_381_reset),
    .io_in(regs_381_io_in),
    .io_init(regs_381_io_init),
    .io_reset(regs_381_io_reset),
    .io_out(regs_381_io_out),
    .io_enable(regs_381_io_enable)
  );
  FF_136 regs_382 (
    .clock(regs_382_clock),
    .reset(regs_382_reset),
    .io_in(regs_382_io_in),
    .io_init(regs_382_io_init),
    .io_reset(regs_382_io_reset),
    .io_out(regs_382_io_out),
    .io_enable(regs_382_io_enable)
  );
  FF_136 regs_383 (
    .clock(regs_383_clock),
    .reset(regs_383_reset),
    .io_in(regs_383_io_in),
    .io_init(regs_383_io_init),
    .io_reset(regs_383_io_reset),
    .io_out(regs_383_io_out),
    .io_enable(regs_383_io_enable)
  );
  FF_136 regs_384 (
    .clock(regs_384_clock),
    .reset(regs_384_reset),
    .io_in(regs_384_io_in),
    .io_init(regs_384_io_init),
    .io_reset(regs_384_io_reset),
    .io_out(regs_384_io_out),
    .io_enable(regs_384_io_enable)
  );
  FF_136 regs_385 (
    .clock(regs_385_clock),
    .reset(regs_385_reset),
    .io_in(regs_385_io_in),
    .io_init(regs_385_io_init),
    .io_reset(regs_385_io_reset),
    .io_out(regs_385_io_out),
    .io_enable(regs_385_io_enable)
  );
  FF_136 regs_386 (
    .clock(regs_386_clock),
    .reset(regs_386_reset),
    .io_in(regs_386_io_in),
    .io_init(regs_386_io_init),
    .io_reset(regs_386_io_reset),
    .io_out(regs_386_io_out),
    .io_enable(regs_386_io_enable)
  );
  FF_136 regs_387 (
    .clock(regs_387_clock),
    .reset(regs_387_reset),
    .io_in(regs_387_io_in),
    .io_init(regs_387_io_init),
    .io_reset(regs_387_io_reset),
    .io_out(regs_387_io_out),
    .io_enable(regs_387_io_enable)
  );
  FF_136 regs_388 (
    .clock(regs_388_clock),
    .reset(regs_388_reset),
    .io_in(regs_388_io_in),
    .io_init(regs_388_io_init),
    .io_reset(regs_388_io_reset),
    .io_out(regs_388_io_out),
    .io_enable(regs_388_io_enable)
  );
  FF_136 regs_389 (
    .clock(regs_389_clock),
    .reset(regs_389_reset),
    .io_in(regs_389_io_in),
    .io_init(regs_389_io_init),
    .io_reset(regs_389_io_reset),
    .io_out(regs_389_io_out),
    .io_enable(regs_389_io_enable)
  );
  FF_136 regs_390 (
    .clock(regs_390_clock),
    .reset(regs_390_reset),
    .io_in(regs_390_io_in),
    .io_init(regs_390_io_init),
    .io_reset(regs_390_io_reset),
    .io_out(regs_390_io_out),
    .io_enable(regs_390_io_enable)
  );
  FF_136 regs_391 (
    .clock(regs_391_clock),
    .reset(regs_391_reset),
    .io_in(regs_391_io_in),
    .io_init(regs_391_io_init),
    .io_reset(regs_391_io_reset),
    .io_out(regs_391_io_out),
    .io_enable(regs_391_io_enable)
  );
  FF_136 regs_392 (
    .clock(regs_392_clock),
    .reset(regs_392_reset),
    .io_in(regs_392_io_in),
    .io_init(regs_392_io_init),
    .io_reset(regs_392_io_reset),
    .io_out(regs_392_io_out),
    .io_enable(regs_392_io_enable)
  );
  FF_136 regs_393 (
    .clock(regs_393_clock),
    .reset(regs_393_reset),
    .io_in(regs_393_io_in),
    .io_init(regs_393_io_init),
    .io_reset(regs_393_io_reset),
    .io_out(regs_393_io_out),
    .io_enable(regs_393_io_enable)
  );
  FF_136 regs_394 (
    .clock(regs_394_clock),
    .reset(regs_394_reset),
    .io_in(regs_394_io_in),
    .io_init(regs_394_io_init),
    .io_reset(regs_394_io_reset),
    .io_out(regs_394_io_out),
    .io_enable(regs_394_io_enable)
  );
  FF_136 regs_395 (
    .clock(regs_395_clock),
    .reset(regs_395_reset),
    .io_in(regs_395_io_in),
    .io_init(regs_395_io_init),
    .io_reset(regs_395_io_reset),
    .io_out(regs_395_io_out),
    .io_enable(regs_395_io_enable)
  );
  FF_136 regs_396 (
    .clock(regs_396_clock),
    .reset(regs_396_reset),
    .io_in(regs_396_io_in),
    .io_init(regs_396_io_init),
    .io_reset(regs_396_io_reset),
    .io_out(regs_396_io_out),
    .io_enable(regs_396_io_enable)
  );
  FF_136 regs_397 (
    .clock(regs_397_clock),
    .reset(regs_397_reset),
    .io_in(regs_397_io_in),
    .io_init(regs_397_io_init),
    .io_reset(regs_397_io_reset),
    .io_out(regs_397_io_out),
    .io_enable(regs_397_io_enable)
  );
  FF_136 regs_398 (
    .clock(regs_398_clock),
    .reset(regs_398_reset),
    .io_in(regs_398_io_in),
    .io_init(regs_398_io_init),
    .io_reset(regs_398_io_reset),
    .io_out(regs_398_io_out),
    .io_enable(regs_398_io_enable)
  );
  FF_136 regs_399 (
    .clock(regs_399_clock),
    .reset(regs_399_reset),
    .io_in(regs_399_io_in),
    .io_init(regs_399_io_init),
    .io_reset(regs_399_io_reset),
    .io_out(regs_399_io_out),
    .io_enable(regs_399_io_enable)
  );
  FF_136 regs_400 (
    .clock(regs_400_clock),
    .reset(regs_400_reset),
    .io_in(regs_400_io_in),
    .io_init(regs_400_io_init),
    .io_reset(regs_400_io_reset),
    .io_out(regs_400_io_out),
    .io_enable(regs_400_io_enable)
  );
  FF_136 regs_401 (
    .clock(regs_401_clock),
    .reset(regs_401_reset),
    .io_in(regs_401_io_in),
    .io_init(regs_401_io_init),
    .io_reset(regs_401_io_reset),
    .io_out(regs_401_io_out),
    .io_enable(regs_401_io_enable)
  );
  FF_136 regs_402 (
    .clock(regs_402_clock),
    .reset(regs_402_reset),
    .io_in(regs_402_io_in),
    .io_init(regs_402_io_init),
    .io_reset(regs_402_io_reset),
    .io_out(regs_402_io_out),
    .io_enable(regs_402_io_enable)
  );
  FF_136 regs_403 (
    .clock(regs_403_clock),
    .reset(regs_403_reset),
    .io_in(regs_403_io_in),
    .io_init(regs_403_io_init),
    .io_reset(regs_403_io_reset),
    .io_out(regs_403_io_out),
    .io_enable(regs_403_io_enable)
  );
  FF_136 regs_404 (
    .clock(regs_404_clock),
    .reset(regs_404_reset),
    .io_in(regs_404_io_in),
    .io_init(regs_404_io_init),
    .io_reset(regs_404_io_reset),
    .io_out(regs_404_io_out),
    .io_enable(regs_404_io_enable)
  );
  FF_136 regs_405 (
    .clock(regs_405_clock),
    .reset(regs_405_reset),
    .io_in(regs_405_io_in),
    .io_init(regs_405_io_init),
    .io_reset(regs_405_io_reset),
    .io_out(regs_405_io_out),
    .io_enable(regs_405_io_enable)
  );
  FF_136 regs_406 (
    .clock(regs_406_clock),
    .reset(regs_406_reset),
    .io_in(regs_406_io_in),
    .io_init(regs_406_io_init),
    .io_reset(regs_406_io_reset),
    .io_out(regs_406_io_out),
    .io_enable(regs_406_io_enable)
  );
  FF_136 regs_407 (
    .clock(regs_407_clock),
    .reset(regs_407_reset),
    .io_in(regs_407_io_in),
    .io_init(regs_407_io_init),
    .io_reset(regs_407_io_reset),
    .io_out(regs_407_io_out),
    .io_enable(regs_407_io_enable)
  );
  FF_136 regs_408 (
    .clock(regs_408_clock),
    .reset(regs_408_reset),
    .io_in(regs_408_io_in),
    .io_init(regs_408_io_init),
    .io_reset(regs_408_io_reset),
    .io_out(regs_408_io_out),
    .io_enable(regs_408_io_enable)
  );
  FF_136 regs_409 (
    .clock(regs_409_clock),
    .reset(regs_409_reset),
    .io_in(regs_409_io_in),
    .io_init(regs_409_io_init),
    .io_reset(regs_409_io_reset),
    .io_out(regs_409_io_out),
    .io_enable(regs_409_io_enable)
  );
  FF_136 regs_410 (
    .clock(regs_410_clock),
    .reset(regs_410_reset),
    .io_in(regs_410_io_in),
    .io_init(regs_410_io_init),
    .io_reset(regs_410_io_reset),
    .io_out(regs_410_io_out),
    .io_enable(regs_410_io_enable)
  );
  FF_136 regs_411 (
    .clock(regs_411_clock),
    .reset(regs_411_reset),
    .io_in(regs_411_io_in),
    .io_init(regs_411_io_init),
    .io_reset(regs_411_io_reset),
    .io_out(regs_411_io_out),
    .io_enable(regs_411_io_enable)
  );
  FF_136 regs_412 (
    .clock(regs_412_clock),
    .reset(regs_412_reset),
    .io_in(regs_412_io_in),
    .io_init(regs_412_io_init),
    .io_reset(regs_412_io_reset),
    .io_out(regs_412_io_out),
    .io_enable(regs_412_io_enable)
  );
  FF_136 regs_413 (
    .clock(regs_413_clock),
    .reset(regs_413_reset),
    .io_in(regs_413_io_in),
    .io_init(regs_413_io_init),
    .io_reset(regs_413_io_reset),
    .io_out(regs_413_io_out),
    .io_enable(regs_413_io_enable)
  );
  FF_136 regs_414 (
    .clock(regs_414_clock),
    .reset(regs_414_reset),
    .io_in(regs_414_io_in),
    .io_init(regs_414_io_init),
    .io_reset(regs_414_io_reset),
    .io_out(regs_414_io_out),
    .io_enable(regs_414_io_enable)
  );
  FF_136 regs_415 (
    .clock(regs_415_clock),
    .reset(regs_415_reset),
    .io_in(regs_415_io_in),
    .io_init(regs_415_io_init),
    .io_reset(regs_415_io_reset),
    .io_out(regs_415_io_out),
    .io_enable(regs_415_io_enable)
  );
  FF_136 regs_416 (
    .clock(regs_416_clock),
    .reset(regs_416_reset),
    .io_in(regs_416_io_in),
    .io_init(regs_416_io_init),
    .io_reset(regs_416_io_reset),
    .io_out(regs_416_io_out),
    .io_enable(regs_416_io_enable)
  );
  FF_136 regs_417 (
    .clock(regs_417_clock),
    .reset(regs_417_reset),
    .io_in(regs_417_io_in),
    .io_init(regs_417_io_init),
    .io_reset(regs_417_io_reset),
    .io_out(regs_417_io_out),
    .io_enable(regs_417_io_enable)
  );
  FF_136 regs_418 (
    .clock(regs_418_clock),
    .reset(regs_418_reset),
    .io_in(regs_418_io_in),
    .io_init(regs_418_io_init),
    .io_reset(regs_418_io_reset),
    .io_out(regs_418_io_out),
    .io_enable(regs_418_io_enable)
  );
  FF_136 regs_419 (
    .clock(regs_419_clock),
    .reset(regs_419_reset),
    .io_in(regs_419_io_in),
    .io_init(regs_419_io_init),
    .io_reset(regs_419_io_reset),
    .io_out(regs_419_io_out),
    .io_enable(regs_419_io_enable)
  );
  FF_136 regs_420 (
    .clock(regs_420_clock),
    .reset(regs_420_reset),
    .io_in(regs_420_io_in),
    .io_init(regs_420_io_init),
    .io_reset(regs_420_io_reset),
    .io_out(regs_420_io_out),
    .io_enable(regs_420_io_enable)
  );
  FF_136 regs_421 (
    .clock(regs_421_clock),
    .reset(regs_421_reset),
    .io_in(regs_421_io_in),
    .io_init(regs_421_io_init),
    .io_reset(regs_421_io_reset),
    .io_out(regs_421_io_out),
    .io_enable(regs_421_io_enable)
  );
  FF_136 regs_422 (
    .clock(regs_422_clock),
    .reset(regs_422_reset),
    .io_in(regs_422_io_in),
    .io_init(regs_422_io_init),
    .io_reset(regs_422_io_reset),
    .io_out(regs_422_io_out),
    .io_enable(regs_422_io_enable)
  );
  FF_136 regs_423 (
    .clock(regs_423_clock),
    .reset(regs_423_reset),
    .io_in(regs_423_io_in),
    .io_init(regs_423_io_init),
    .io_reset(regs_423_io_reset),
    .io_out(regs_423_io_out),
    .io_enable(regs_423_io_enable)
  );
  FF_136 regs_424 (
    .clock(regs_424_clock),
    .reset(regs_424_reset),
    .io_in(regs_424_io_in),
    .io_init(regs_424_io_init),
    .io_reset(regs_424_io_reset),
    .io_out(regs_424_io_out),
    .io_enable(regs_424_io_enable)
  );
  FF_136 regs_425 (
    .clock(regs_425_clock),
    .reset(regs_425_reset),
    .io_in(regs_425_io_in),
    .io_init(regs_425_io_init),
    .io_reset(regs_425_io_reset),
    .io_out(regs_425_io_out),
    .io_enable(regs_425_io_enable)
  );
  FF_136 regs_426 (
    .clock(regs_426_clock),
    .reset(regs_426_reset),
    .io_in(regs_426_io_in),
    .io_init(regs_426_io_init),
    .io_reset(regs_426_io_reset),
    .io_out(regs_426_io_out),
    .io_enable(regs_426_io_enable)
  );
  FF_136 regs_427 (
    .clock(regs_427_clock),
    .reset(regs_427_reset),
    .io_in(regs_427_io_in),
    .io_init(regs_427_io_init),
    .io_reset(regs_427_io_reset),
    .io_out(regs_427_io_out),
    .io_enable(regs_427_io_enable)
  );
  FF_136 regs_428 (
    .clock(regs_428_clock),
    .reset(regs_428_reset),
    .io_in(regs_428_io_in),
    .io_init(regs_428_io_init),
    .io_reset(regs_428_io_reset),
    .io_out(regs_428_io_out),
    .io_enable(regs_428_io_enable)
  );
  FF_136 regs_429 (
    .clock(regs_429_clock),
    .reset(regs_429_reset),
    .io_in(regs_429_io_in),
    .io_init(regs_429_io_init),
    .io_reset(regs_429_io_reset),
    .io_out(regs_429_io_out),
    .io_enable(regs_429_io_enable)
  );
  FF_136 regs_430 (
    .clock(regs_430_clock),
    .reset(regs_430_reset),
    .io_in(regs_430_io_in),
    .io_init(regs_430_io_init),
    .io_reset(regs_430_io_reset),
    .io_out(regs_430_io_out),
    .io_enable(regs_430_io_enable)
  );
  FF_136 regs_431 (
    .clock(regs_431_clock),
    .reset(regs_431_reset),
    .io_in(regs_431_io_in),
    .io_init(regs_431_io_init),
    .io_reset(regs_431_io_reset),
    .io_out(regs_431_io_out),
    .io_enable(regs_431_io_enable)
  );
  FF_136 regs_432 (
    .clock(regs_432_clock),
    .reset(regs_432_reset),
    .io_in(regs_432_io_in),
    .io_init(regs_432_io_init),
    .io_reset(regs_432_io_reset),
    .io_out(regs_432_io_out),
    .io_enable(regs_432_io_enable)
  );
  FF_136 regs_433 (
    .clock(regs_433_clock),
    .reset(regs_433_reset),
    .io_in(regs_433_io_in),
    .io_init(regs_433_io_init),
    .io_reset(regs_433_io_reset),
    .io_out(regs_433_io_out),
    .io_enable(regs_433_io_enable)
  );
  FF_136 regs_434 (
    .clock(regs_434_clock),
    .reset(regs_434_reset),
    .io_in(regs_434_io_in),
    .io_init(regs_434_io_init),
    .io_reset(regs_434_io_reset),
    .io_out(regs_434_io_out),
    .io_enable(regs_434_io_enable)
  );
  FF_136 regs_435 (
    .clock(regs_435_clock),
    .reset(regs_435_reset),
    .io_in(regs_435_io_in),
    .io_init(regs_435_io_init),
    .io_reset(regs_435_io_reset),
    .io_out(regs_435_io_out),
    .io_enable(regs_435_io_enable)
  );
  FF_136 regs_436 (
    .clock(regs_436_clock),
    .reset(regs_436_reset),
    .io_in(regs_436_io_in),
    .io_init(regs_436_io_init),
    .io_reset(regs_436_io_reset),
    .io_out(regs_436_io_out),
    .io_enable(regs_436_io_enable)
  );
  FF_136 regs_437 (
    .clock(regs_437_clock),
    .reset(regs_437_reset),
    .io_in(regs_437_io_in),
    .io_init(regs_437_io_init),
    .io_reset(regs_437_io_reset),
    .io_out(regs_437_io_out),
    .io_enable(regs_437_io_enable)
  );
  FF_136 regs_438 (
    .clock(regs_438_clock),
    .reset(regs_438_reset),
    .io_in(regs_438_io_in),
    .io_init(regs_438_io_init),
    .io_reset(regs_438_io_reset),
    .io_out(regs_438_io_out),
    .io_enable(regs_438_io_enable)
  );
  FF_136 regs_439 (
    .clock(regs_439_clock),
    .reset(regs_439_reset),
    .io_in(regs_439_io_in),
    .io_init(regs_439_io_init),
    .io_reset(regs_439_io_reset),
    .io_out(regs_439_io_out),
    .io_enable(regs_439_io_enable)
  );
  FF_136 regs_440 (
    .clock(regs_440_clock),
    .reset(regs_440_reset),
    .io_in(regs_440_io_in),
    .io_init(regs_440_io_init),
    .io_reset(regs_440_io_reset),
    .io_out(regs_440_io_out),
    .io_enable(regs_440_io_enable)
  );
  FF_136 regs_441 (
    .clock(regs_441_clock),
    .reset(regs_441_reset),
    .io_in(regs_441_io_in),
    .io_init(regs_441_io_init),
    .io_reset(regs_441_io_reset),
    .io_out(regs_441_io_out),
    .io_enable(regs_441_io_enable)
  );
  FF_136 regs_442 (
    .clock(regs_442_clock),
    .reset(regs_442_reset),
    .io_in(regs_442_io_in),
    .io_init(regs_442_io_init),
    .io_reset(regs_442_io_reset),
    .io_out(regs_442_io_out),
    .io_enable(regs_442_io_enable)
  );
  FF_136 regs_443 (
    .clock(regs_443_clock),
    .reset(regs_443_reset),
    .io_in(regs_443_io_in),
    .io_init(regs_443_io_init),
    .io_reset(regs_443_io_reset),
    .io_out(regs_443_io_out),
    .io_enable(regs_443_io_enable)
  );
  FF_136 regs_444 (
    .clock(regs_444_clock),
    .reset(regs_444_reset),
    .io_in(regs_444_io_in),
    .io_init(regs_444_io_init),
    .io_reset(regs_444_io_reset),
    .io_out(regs_444_io_out),
    .io_enable(regs_444_io_enable)
  );
  FF_136 regs_445 (
    .clock(regs_445_clock),
    .reset(regs_445_reset),
    .io_in(regs_445_io_in),
    .io_init(regs_445_io_init),
    .io_reset(regs_445_io_reset),
    .io_out(regs_445_io_out),
    .io_enable(regs_445_io_enable)
  );
  FF_136 regs_446 (
    .clock(regs_446_clock),
    .reset(regs_446_reset),
    .io_in(regs_446_io_in),
    .io_init(regs_446_io_init),
    .io_reset(regs_446_io_reset),
    .io_out(regs_446_io_out),
    .io_enable(regs_446_io_enable)
  );
  FF_136 regs_447 (
    .clock(regs_447_clock),
    .reset(regs_447_reset),
    .io_in(regs_447_io_in),
    .io_init(regs_447_io_init),
    .io_reset(regs_447_io_reset),
    .io_out(regs_447_io_out),
    .io_enable(regs_447_io_enable)
  );
  FF_136 regs_448 (
    .clock(regs_448_clock),
    .reset(regs_448_reset),
    .io_in(regs_448_io_in),
    .io_init(regs_448_io_init),
    .io_reset(regs_448_io_reset),
    .io_out(regs_448_io_out),
    .io_enable(regs_448_io_enable)
  );
  FF_136 regs_449 (
    .clock(regs_449_clock),
    .reset(regs_449_reset),
    .io_in(regs_449_io_in),
    .io_init(regs_449_io_init),
    .io_reset(regs_449_io_reset),
    .io_out(regs_449_io_out),
    .io_enable(regs_449_io_enable)
  );
  FF_136 regs_450 (
    .clock(regs_450_clock),
    .reset(regs_450_reset),
    .io_in(regs_450_io_in),
    .io_init(regs_450_io_init),
    .io_reset(regs_450_io_reset),
    .io_out(regs_450_io_out),
    .io_enable(regs_450_io_enable)
  );
  FF_136 regs_451 (
    .clock(regs_451_clock),
    .reset(regs_451_reset),
    .io_in(regs_451_io_in),
    .io_init(regs_451_io_init),
    .io_reset(regs_451_io_reset),
    .io_out(regs_451_io_out),
    .io_enable(regs_451_io_enable)
  );
  FF_136 regs_452 (
    .clock(regs_452_clock),
    .reset(regs_452_reset),
    .io_in(regs_452_io_in),
    .io_init(regs_452_io_init),
    .io_reset(regs_452_io_reset),
    .io_out(regs_452_io_out),
    .io_enable(regs_452_io_enable)
  );
  FF_136 regs_453 (
    .clock(regs_453_clock),
    .reset(regs_453_reset),
    .io_in(regs_453_io_in),
    .io_init(regs_453_io_init),
    .io_reset(regs_453_io_reset),
    .io_out(regs_453_io_out),
    .io_enable(regs_453_io_enable)
  );
  FF_136 regs_454 (
    .clock(regs_454_clock),
    .reset(regs_454_reset),
    .io_in(regs_454_io_in),
    .io_init(regs_454_io_init),
    .io_reset(regs_454_io_reset),
    .io_out(regs_454_io_out),
    .io_enable(regs_454_io_enable)
  );
  FF_136 regs_455 (
    .clock(regs_455_clock),
    .reset(regs_455_reset),
    .io_in(regs_455_io_in),
    .io_init(regs_455_io_init),
    .io_reset(regs_455_io_reset),
    .io_out(regs_455_io_out),
    .io_enable(regs_455_io_enable)
  );
  FF_136 regs_456 (
    .clock(regs_456_clock),
    .reset(regs_456_reset),
    .io_in(regs_456_io_in),
    .io_init(regs_456_io_init),
    .io_reset(regs_456_io_reset),
    .io_out(regs_456_io_out),
    .io_enable(regs_456_io_enable)
  );
  FF_136 regs_457 (
    .clock(regs_457_clock),
    .reset(regs_457_reset),
    .io_in(regs_457_io_in),
    .io_init(regs_457_io_init),
    .io_reset(regs_457_io_reset),
    .io_out(regs_457_io_out),
    .io_enable(regs_457_io_enable)
  );
  FF_136 regs_458 (
    .clock(regs_458_clock),
    .reset(regs_458_reset),
    .io_in(regs_458_io_in),
    .io_init(regs_458_io_init),
    .io_reset(regs_458_io_reset),
    .io_out(regs_458_io_out),
    .io_enable(regs_458_io_enable)
  );
  FF_136 regs_459 (
    .clock(regs_459_clock),
    .reset(regs_459_reset),
    .io_in(regs_459_io_in),
    .io_init(regs_459_io_init),
    .io_reset(regs_459_io_reset),
    .io_out(regs_459_io_out),
    .io_enable(regs_459_io_enable)
  );
  FF_136 regs_460 (
    .clock(regs_460_clock),
    .reset(regs_460_reset),
    .io_in(regs_460_io_in),
    .io_init(regs_460_io_init),
    .io_reset(regs_460_io_reset),
    .io_out(regs_460_io_out),
    .io_enable(regs_460_io_enable)
  );
  FF_136 regs_461 (
    .clock(regs_461_clock),
    .reset(regs_461_reset),
    .io_in(regs_461_io_in),
    .io_init(regs_461_io_init),
    .io_reset(regs_461_io_reset),
    .io_out(regs_461_io_out),
    .io_enable(regs_461_io_enable)
  );
  FF_136 regs_462 (
    .clock(regs_462_clock),
    .reset(regs_462_reset),
    .io_in(regs_462_io_in),
    .io_init(regs_462_io_init),
    .io_reset(regs_462_io_reset),
    .io_out(regs_462_io_out),
    .io_enable(regs_462_io_enable)
  );
  FF_136 regs_463 (
    .clock(regs_463_clock),
    .reset(regs_463_reset),
    .io_in(regs_463_io_in),
    .io_init(regs_463_io_init),
    .io_reset(regs_463_io_reset),
    .io_out(regs_463_io_out),
    .io_enable(regs_463_io_enable)
  );
  FF_136 regs_464 (
    .clock(regs_464_clock),
    .reset(regs_464_reset),
    .io_in(regs_464_io_in),
    .io_init(regs_464_io_init),
    .io_reset(regs_464_io_reset),
    .io_out(regs_464_io_out),
    .io_enable(regs_464_io_enable)
  );
  FF_136 regs_465 (
    .clock(regs_465_clock),
    .reset(regs_465_reset),
    .io_in(regs_465_io_in),
    .io_init(regs_465_io_init),
    .io_reset(regs_465_io_reset),
    .io_out(regs_465_io_out),
    .io_enable(regs_465_io_enable)
  );
  FF_136 regs_466 (
    .clock(regs_466_clock),
    .reset(regs_466_reset),
    .io_in(regs_466_io_in),
    .io_init(regs_466_io_init),
    .io_reset(regs_466_io_reset),
    .io_out(regs_466_io_out),
    .io_enable(regs_466_io_enable)
  );
  FF_136 regs_467 (
    .clock(regs_467_clock),
    .reset(regs_467_reset),
    .io_in(regs_467_io_in),
    .io_init(regs_467_io_init),
    .io_reset(regs_467_io_reset),
    .io_out(regs_467_io_out),
    .io_enable(regs_467_io_enable)
  );
  FF_136 regs_468 (
    .clock(regs_468_clock),
    .reset(regs_468_reset),
    .io_in(regs_468_io_in),
    .io_init(regs_468_io_init),
    .io_reset(regs_468_io_reset),
    .io_out(regs_468_io_out),
    .io_enable(regs_468_io_enable)
  );
  FF_136 regs_469 (
    .clock(regs_469_clock),
    .reset(regs_469_reset),
    .io_in(regs_469_io_in),
    .io_init(regs_469_io_init),
    .io_reset(regs_469_io_reset),
    .io_out(regs_469_io_out),
    .io_enable(regs_469_io_enable)
  );
  FF_136 regs_470 (
    .clock(regs_470_clock),
    .reset(regs_470_reset),
    .io_in(regs_470_io_in),
    .io_init(regs_470_io_init),
    .io_reset(regs_470_io_reset),
    .io_out(regs_470_io_out),
    .io_enable(regs_470_io_enable)
  );
  FF_136 regs_471 (
    .clock(regs_471_clock),
    .reset(regs_471_reset),
    .io_in(regs_471_io_in),
    .io_init(regs_471_io_init),
    .io_reset(regs_471_io_reset),
    .io_out(regs_471_io_out),
    .io_enable(regs_471_io_enable)
  );
  FF_136 regs_472 (
    .clock(regs_472_clock),
    .reset(regs_472_reset),
    .io_in(regs_472_io_in),
    .io_init(regs_472_io_init),
    .io_reset(regs_472_io_reset),
    .io_out(regs_472_io_out),
    .io_enable(regs_472_io_enable)
  );
  FF_136 regs_473 (
    .clock(regs_473_clock),
    .reset(regs_473_reset),
    .io_in(regs_473_io_in),
    .io_init(regs_473_io_init),
    .io_reset(regs_473_io_reset),
    .io_out(regs_473_io_out),
    .io_enable(regs_473_io_enable)
  );
  FF_136 regs_474 (
    .clock(regs_474_clock),
    .reset(regs_474_reset),
    .io_in(regs_474_io_in),
    .io_init(regs_474_io_init),
    .io_reset(regs_474_io_reset),
    .io_out(regs_474_io_out),
    .io_enable(regs_474_io_enable)
  );
  FF_136 regs_475 (
    .clock(regs_475_clock),
    .reset(regs_475_reset),
    .io_in(regs_475_io_in),
    .io_init(regs_475_io_init),
    .io_reset(regs_475_io_reset),
    .io_out(regs_475_io_out),
    .io_enable(regs_475_io_enable)
  );
  FF_136 regs_476 (
    .clock(regs_476_clock),
    .reset(regs_476_reset),
    .io_in(regs_476_io_in),
    .io_init(regs_476_io_init),
    .io_reset(regs_476_io_reset),
    .io_out(regs_476_io_out),
    .io_enable(regs_476_io_enable)
  );
  FF_136 regs_477 (
    .clock(regs_477_clock),
    .reset(regs_477_reset),
    .io_in(regs_477_io_in),
    .io_init(regs_477_io_init),
    .io_reset(regs_477_io_reset),
    .io_out(regs_477_io_out),
    .io_enable(regs_477_io_enable)
  );
  FF_136 regs_478 (
    .clock(regs_478_clock),
    .reset(regs_478_reset),
    .io_in(regs_478_io_in),
    .io_init(regs_478_io_init),
    .io_reset(regs_478_io_reset),
    .io_out(regs_478_io_out),
    .io_enable(regs_478_io_enable)
  );
  FF_136 regs_479 (
    .clock(regs_479_clock),
    .reset(regs_479_reset),
    .io_in(regs_479_io_in),
    .io_init(regs_479_io_init),
    .io_reset(regs_479_io_reset),
    .io_out(regs_479_io_out),
    .io_enable(regs_479_io_enable)
  );
  FF_136 regs_480 (
    .clock(regs_480_clock),
    .reset(regs_480_reset),
    .io_in(regs_480_io_in),
    .io_init(regs_480_io_init),
    .io_reset(regs_480_io_reset),
    .io_out(regs_480_io_out),
    .io_enable(regs_480_io_enable)
  );
  FF_136 regs_481 (
    .clock(regs_481_clock),
    .reset(regs_481_reset),
    .io_in(regs_481_io_in),
    .io_init(regs_481_io_init),
    .io_reset(regs_481_io_reset),
    .io_out(regs_481_io_out),
    .io_enable(regs_481_io_enable)
  );
  FF_136 regs_482 (
    .clock(regs_482_clock),
    .reset(regs_482_reset),
    .io_in(regs_482_io_in),
    .io_init(regs_482_io_init),
    .io_reset(regs_482_io_reset),
    .io_out(regs_482_io_out),
    .io_enable(regs_482_io_enable)
  );
  FF_136 regs_483 (
    .clock(regs_483_clock),
    .reset(regs_483_reset),
    .io_in(regs_483_io_in),
    .io_init(regs_483_io_init),
    .io_reset(regs_483_io_reset),
    .io_out(regs_483_io_out),
    .io_enable(regs_483_io_enable)
  );
  FF_136 regs_484 (
    .clock(regs_484_clock),
    .reset(regs_484_reset),
    .io_in(regs_484_io_in),
    .io_init(regs_484_io_init),
    .io_reset(regs_484_io_reset),
    .io_out(regs_484_io_out),
    .io_enable(regs_484_io_enable)
  );
  FF_136 regs_485 (
    .clock(regs_485_clock),
    .reset(regs_485_reset),
    .io_in(regs_485_io_in),
    .io_init(regs_485_io_init),
    .io_reset(regs_485_io_reset),
    .io_out(regs_485_io_out),
    .io_enable(regs_485_io_enable)
  );
  FF_136 regs_486 (
    .clock(regs_486_clock),
    .reset(regs_486_reset),
    .io_in(regs_486_io_in),
    .io_init(regs_486_io_init),
    .io_reset(regs_486_io_reset),
    .io_out(regs_486_io_out),
    .io_enable(regs_486_io_enable)
  );
  FF_136 regs_487 (
    .clock(regs_487_clock),
    .reset(regs_487_reset),
    .io_in(regs_487_io_in),
    .io_init(regs_487_io_init),
    .io_reset(regs_487_io_reset),
    .io_out(regs_487_io_out),
    .io_enable(regs_487_io_enable)
  );
  FF_136 regs_488 (
    .clock(regs_488_clock),
    .reset(regs_488_reset),
    .io_in(regs_488_io_in),
    .io_init(regs_488_io_init),
    .io_reset(regs_488_io_reset),
    .io_out(regs_488_io_out),
    .io_enable(regs_488_io_enable)
  );
  FF_136 regs_489 (
    .clock(regs_489_clock),
    .reset(regs_489_reset),
    .io_in(regs_489_io_in),
    .io_init(regs_489_io_init),
    .io_reset(regs_489_io_reset),
    .io_out(regs_489_io_out),
    .io_enable(regs_489_io_enable)
  );
  FF_136 regs_490 (
    .clock(regs_490_clock),
    .reset(regs_490_reset),
    .io_in(regs_490_io_in),
    .io_init(regs_490_io_init),
    .io_reset(regs_490_io_reset),
    .io_out(regs_490_io_out),
    .io_enable(regs_490_io_enable)
  );
  FF_136 regs_491 (
    .clock(regs_491_clock),
    .reset(regs_491_reset),
    .io_in(regs_491_io_in),
    .io_init(regs_491_io_init),
    .io_reset(regs_491_io_reset),
    .io_out(regs_491_io_out),
    .io_enable(regs_491_io_enable)
  );
  FF_136 regs_492 (
    .clock(regs_492_clock),
    .reset(regs_492_reset),
    .io_in(regs_492_io_in),
    .io_init(regs_492_io_init),
    .io_reset(regs_492_io_reset),
    .io_out(regs_492_io_out),
    .io_enable(regs_492_io_enable)
  );
  FF_136 regs_493 (
    .clock(regs_493_clock),
    .reset(regs_493_reset),
    .io_in(regs_493_io_in),
    .io_init(regs_493_io_init),
    .io_reset(regs_493_io_reset),
    .io_out(regs_493_io_out),
    .io_enable(regs_493_io_enable)
  );
  FF_136 regs_494 (
    .clock(regs_494_clock),
    .reset(regs_494_reset),
    .io_in(regs_494_io_in),
    .io_init(regs_494_io_init),
    .io_reset(regs_494_io_reset),
    .io_out(regs_494_io_out),
    .io_enable(regs_494_io_enable)
  );
  FF_136 regs_495 (
    .clock(regs_495_clock),
    .reset(regs_495_reset),
    .io_in(regs_495_io_in),
    .io_init(regs_495_io_init),
    .io_reset(regs_495_io_reset),
    .io_out(regs_495_io_out),
    .io_enable(regs_495_io_enable)
  );
  FF_136 regs_496 (
    .clock(regs_496_clock),
    .reset(regs_496_reset),
    .io_in(regs_496_io_in),
    .io_init(regs_496_io_init),
    .io_reset(regs_496_io_reset),
    .io_out(regs_496_io_out),
    .io_enable(regs_496_io_enable)
  );
  FF_136 regs_497 (
    .clock(regs_497_clock),
    .reset(regs_497_reset),
    .io_in(regs_497_io_in),
    .io_init(regs_497_io_init),
    .io_reset(regs_497_io_reset),
    .io_out(regs_497_io_out),
    .io_enable(regs_497_io_enable)
  );
  FF_136 regs_498 (
    .clock(regs_498_clock),
    .reset(regs_498_reset),
    .io_in(regs_498_io_in),
    .io_init(regs_498_io_init),
    .io_reset(regs_498_io_reset),
    .io_out(regs_498_io_out),
    .io_enable(regs_498_io_enable)
  );
  FF_136 regs_499 (
    .clock(regs_499_clock),
    .reset(regs_499_reset),
    .io_in(regs_499_io_in),
    .io_init(regs_499_io_init),
    .io_reset(regs_499_io_reset),
    .io_out(regs_499_io_out),
    .io_enable(regs_499_io_enable)
  );
  FF_136 regs_500 (
    .clock(regs_500_clock),
    .reset(regs_500_reset),
    .io_in(regs_500_io_in),
    .io_init(regs_500_io_init),
    .io_reset(regs_500_io_reset),
    .io_out(regs_500_io_out),
    .io_enable(regs_500_io_enable)
  );
  FF_136 regs_501 (
    .clock(regs_501_clock),
    .reset(regs_501_reset),
    .io_in(regs_501_io_in),
    .io_init(regs_501_io_init),
    .io_reset(regs_501_io_reset),
    .io_out(regs_501_io_out),
    .io_enable(regs_501_io_enable)
  );
  FF_136 regs_502 (
    .clock(regs_502_clock),
    .reset(regs_502_reset),
    .io_in(regs_502_io_in),
    .io_init(regs_502_io_init),
    .io_reset(regs_502_io_reset),
    .io_out(regs_502_io_out),
    .io_enable(regs_502_io_enable)
  );
  FF_136 regs_503 (
    .clock(regs_503_clock),
    .reset(regs_503_reset),
    .io_in(regs_503_io_in),
    .io_init(regs_503_io_init),
    .io_reset(regs_503_io_reset),
    .io_out(regs_503_io_out),
    .io_enable(regs_503_io_enable)
  );
  FF_136 regs_504 (
    .clock(regs_504_clock),
    .reset(regs_504_reset),
    .io_in(regs_504_io_in),
    .io_init(regs_504_io_init),
    .io_reset(regs_504_io_reset),
    .io_out(regs_504_io_out),
    .io_enable(regs_504_io_enable)
  );
  FF_136 regs_505 (
    .clock(regs_505_clock),
    .reset(regs_505_reset),
    .io_in(regs_505_io_in),
    .io_init(regs_505_io_init),
    .io_reset(regs_505_io_reset),
    .io_out(regs_505_io_out),
    .io_enable(regs_505_io_enable)
  );
  MuxN_80 rport (
    .io_ins_0(rport_io_ins_0),
    .io_ins_1(rport_io_ins_1),
    .io_ins_2(rport_io_ins_2),
    .io_ins_3(rport_io_ins_3),
    .io_ins_4(rport_io_ins_4),
    .io_ins_5(rport_io_ins_5),
    .io_ins_6(rport_io_ins_6),
    .io_ins_7(rport_io_ins_7),
    .io_ins_8(rport_io_ins_8),
    .io_ins_9(rport_io_ins_9),
    .io_ins_10(rport_io_ins_10),
    .io_ins_11(rport_io_ins_11),
    .io_ins_12(rport_io_ins_12),
    .io_ins_13(rport_io_ins_13),
    .io_ins_14(rport_io_ins_14),
    .io_ins_15(rport_io_ins_15),
    .io_ins_16(rport_io_ins_16),
    .io_ins_17(rport_io_ins_17),
    .io_ins_18(rport_io_ins_18),
    .io_ins_19(rport_io_ins_19),
    .io_ins_20(rport_io_ins_20),
    .io_ins_21(rport_io_ins_21),
    .io_ins_22(rport_io_ins_22),
    .io_ins_23(rport_io_ins_23),
    .io_ins_24(rport_io_ins_24),
    .io_ins_25(rport_io_ins_25),
    .io_ins_26(rport_io_ins_26),
    .io_ins_27(rport_io_ins_27),
    .io_ins_28(rport_io_ins_28),
    .io_ins_29(rport_io_ins_29),
    .io_ins_30(rport_io_ins_30),
    .io_ins_31(rport_io_ins_31),
    .io_ins_32(rport_io_ins_32),
    .io_ins_33(rport_io_ins_33),
    .io_ins_34(rport_io_ins_34),
    .io_ins_35(rport_io_ins_35),
    .io_ins_36(rport_io_ins_36),
    .io_ins_37(rport_io_ins_37),
    .io_ins_38(rport_io_ins_38),
    .io_ins_39(rport_io_ins_39),
    .io_ins_40(rport_io_ins_40),
    .io_ins_41(rport_io_ins_41),
    .io_ins_42(rport_io_ins_42),
    .io_ins_43(rport_io_ins_43),
    .io_ins_44(rport_io_ins_44),
    .io_ins_45(rport_io_ins_45),
    .io_ins_46(rport_io_ins_46),
    .io_ins_47(rport_io_ins_47),
    .io_ins_48(rport_io_ins_48),
    .io_ins_49(rport_io_ins_49),
    .io_ins_50(rport_io_ins_50),
    .io_ins_51(rport_io_ins_51),
    .io_ins_52(rport_io_ins_52),
    .io_ins_53(rport_io_ins_53),
    .io_ins_54(rport_io_ins_54),
    .io_ins_55(rport_io_ins_55),
    .io_ins_56(rport_io_ins_56),
    .io_ins_57(rport_io_ins_57),
    .io_ins_58(rport_io_ins_58),
    .io_ins_59(rport_io_ins_59),
    .io_ins_60(rport_io_ins_60),
    .io_ins_61(rport_io_ins_61),
    .io_ins_62(rport_io_ins_62),
    .io_ins_63(rport_io_ins_63),
    .io_ins_64(rport_io_ins_64),
    .io_ins_65(rport_io_ins_65),
    .io_ins_66(rport_io_ins_66),
    .io_ins_67(rport_io_ins_67),
    .io_ins_68(rport_io_ins_68),
    .io_ins_69(rport_io_ins_69),
    .io_ins_70(rport_io_ins_70),
    .io_ins_71(rport_io_ins_71),
    .io_ins_72(rport_io_ins_72),
    .io_ins_73(rport_io_ins_73),
    .io_ins_74(rport_io_ins_74),
    .io_ins_75(rport_io_ins_75),
    .io_ins_76(rport_io_ins_76),
    .io_ins_77(rport_io_ins_77),
    .io_ins_78(rport_io_ins_78),
    .io_ins_79(rport_io_ins_79),
    .io_ins_80(rport_io_ins_80),
    .io_ins_81(rport_io_ins_81),
    .io_ins_82(rport_io_ins_82),
    .io_ins_83(rport_io_ins_83),
    .io_ins_84(rport_io_ins_84),
    .io_ins_85(rport_io_ins_85),
    .io_ins_86(rport_io_ins_86),
    .io_ins_87(rport_io_ins_87),
    .io_ins_88(rport_io_ins_88),
    .io_ins_89(rport_io_ins_89),
    .io_ins_90(rport_io_ins_90),
    .io_ins_91(rport_io_ins_91),
    .io_ins_92(rport_io_ins_92),
    .io_ins_93(rport_io_ins_93),
    .io_ins_94(rport_io_ins_94),
    .io_ins_95(rport_io_ins_95),
    .io_ins_96(rport_io_ins_96),
    .io_ins_97(rport_io_ins_97),
    .io_ins_98(rport_io_ins_98),
    .io_ins_99(rport_io_ins_99),
    .io_ins_100(rport_io_ins_100),
    .io_ins_101(rport_io_ins_101),
    .io_ins_102(rport_io_ins_102),
    .io_ins_103(rport_io_ins_103),
    .io_ins_104(rport_io_ins_104),
    .io_ins_105(rport_io_ins_105),
    .io_ins_106(rport_io_ins_106),
    .io_ins_107(rport_io_ins_107),
    .io_ins_108(rport_io_ins_108),
    .io_ins_109(rport_io_ins_109),
    .io_ins_110(rport_io_ins_110),
    .io_ins_111(rport_io_ins_111),
    .io_ins_112(rport_io_ins_112),
    .io_ins_113(rport_io_ins_113),
    .io_ins_114(rport_io_ins_114),
    .io_ins_115(rport_io_ins_115),
    .io_ins_116(rport_io_ins_116),
    .io_ins_117(rport_io_ins_117),
    .io_ins_118(rport_io_ins_118),
    .io_ins_119(rport_io_ins_119),
    .io_ins_120(rport_io_ins_120),
    .io_ins_121(rport_io_ins_121),
    .io_ins_122(rport_io_ins_122),
    .io_ins_123(rport_io_ins_123),
    .io_ins_124(rport_io_ins_124),
    .io_ins_125(rport_io_ins_125),
    .io_ins_126(rport_io_ins_126),
    .io_ins_127(rport_io_ins_127),
    .io_ins_128(rport_io_ins_128),
    .io_ins_129(rport_io_ins_129),
    .io_ins_130(rport_io_ins_130),
    .io_ins_131(rport_io_ins_131),
    .io_ins_132(rport_io_ins_132),
    .io_ins_133(rport_io_ins_133),
    .io_ins_134(rport_io_ins_134),
    .io_ins_135(rport_io_ins_135),
    .io_ins_136(rport_io_ins_136),
    .io_ins_137(rport_io_ins_137),
    .io_ins_138(rport_io_ins_138),
    .io_ins_139(rport_io_ins_139),
    .io_ins_140(rport_io_ins_140),
    .io_ins_141(rport_io_ins_141),
    .io_ins_142(rport_io_ins_142),
    .io_ins_143(rport_io_ins_143),
    .io_ins_144(rport_io_ins_144),
    .io_ins_145(rport_io_ins_145),
    .io_ins_146(rport_io_ins_146),
    .io_ins_147(rport_io_ins_147),
    .io_ins_148(rport_io_ins_148),
    .io_ins_149(rport_io_ins_149),
    .io_ins_150(rport_io_ins_150),
    .io_ins_151(rport_io_ins_151),
    .io_ins_152(rport_io_ins_152),
    .io_ins_153(rport_io_ins_153),
    .io_ins_154(rport_io_ins_154),
    .io_ins_155(rport_io_ins_155),
    .io_ins_156(rport_io_ins_156),
    .io_ins_157(rport_io_ins_157),
    .io_ins_158(rport_io_ins_158),
    .io_ins_159(rport_io_ins_159),
    .io_ins_160(rport_io_ins_160),
    .io_ins_161(rport_io_ins_161),
    .io_ins_162(rport_io_ins_162),
    .io_ins_163(rport_io_ins_163),
    .io_ins_164(rport_io_ins_164),
    .io_ins_165(rport_io_ins_165),
    .io_ins_166(rport_io_ins_166),
    .io_ins_167(rport_io_ins_167),
    .io_ins_168(rport_io_ins_168),
    .io_ins_169(rport_io_ins_169),
    .io_ins_170(rport_io_ins_170),
    .io_ins_171(rport_io_ins_171),
    .io_ins_172(rport_io_ins_172),
    .io_ins_173(rport_io_ins_173),
    .io_ins_174(rport_io_ins_174),
    .io_ins_175(rport_io_ins_175),
    .io_ins_176(rport_io_ins_176),
    .io_ins_177(rport_io_ins_177),
    .io_ins_178(rport_io_ins_178),
    .io_ins_179(rport_io_ins_179),
    .io_ins_180(rport_io_ins_180),
    .io_ins_181(rport_io_ins_181),
    .io_ins_182(rport_io_ins_182),
    .io_ins_183(rport_io_ins_183),
    .io_ins_184(rport_io_ins_184),
    .io_ins_185(rport_io_ins_185),
    .io_ins_186(rport_io_ins_186),
    .io_ins_187(rport_io_ins_187),
    .io_ins_188(rport_io_ins_188),
    .io_ins_189(rport_io_ins_189),
    .io_ins_190(rport_io_ins_190),
    .io_ins_191(rport_io_ins_191),
    .io_ins_192(rport_io_ins_192),
    .io_ins_193(rport_io_ins_193),
    .io_ins_194(rport_io_ins_194),
    .io_ins_195(rport_io_ins_195),
    .io_ins_196(rport_io_ins_196),
    .io_ins_197(rport_io_ins_197),
    .io_ins_198(rport_io_ins_198),
    .io_ins_199(rport_io_ins_199),
    .io_ins_200(rport_io_ins_200),
    .io_ins_201(rport_io_ins_201),
    .io_ins_202(rport_io_ins_202),
    .io_ins_203(rport_io_ins_203),
    .io_ins_204(rport_io_ins_204),
    .io_ins_205(rport_io_ins_205),
    .io_ins_206(rport_io_ins_206),
    .io_ins_207(rport_io_ins_207),
    .io_ins_208(rport_io_ins_208),
    .io_ins_209(rport_io_ins_209),
    .io_ins_210(rport_io_ins_210),
    .io_ins_211(rport_io_ins_211),
    .io_ins_212(rport_io_ins_212),
    .io_ins_213(rport_io_ins_213),
    .io_ins_214(rport_io_ins_214),
    .io_ins_215(rport_io_ins_215),
    .io_ins_216(rport_io_ins_216),
    .io_ins_217(rport_io_ins_217),
    .io_ins_218(rport_io_ins_218),
    .io_ins_219(rport_io_ins_219),
    .io_ins_220(rport_io_ins_220),
    .io_ins_221(rport_io_ins_221),
    .io_ins_222(rport_io_ins_222),
    .io_ins_223(rport_io_ins_223),
    .io_ins_224(rport_io_ins_224),
    .io_ins_225(rport_io_ins_225),
    .io_ins_226(rport_io_ins_226),
    .io_ins_227(rport_io_ins_227),
    .io_ins_228(rport_io_ins_228),
    .io_ins_229(rport_io_ins_229),
    .io_ins_230(rport_io_ins_230),
    .io_ins_231(rport_io_ins_231),
    .io_ins_232(rport_io_ins_232),
    .io_ins_233(rport_io_ins_233),
    .io_ins_234(rport_io_ins_234),
    .io_ins_235(rport_io_ins_235),
    .io_ins_236(rport_io_ins_236),
    .io_ins_237(rport_io_ins_237),
    .io_ins_238(rport_io_ins_238),
    .io_ins_239(rport_io_ins_239),
    .io_ins_240(rport_io_ins_240),
    .io_ins_241(rport_io_ins_241),
    .io_ins_242(rport_io_ins_242),
    .io_ins_243(rport_io_ins_243),
    .io_ins_244(rport_io_ins_244),
    .io_ins_245(rport_io_ins_245),
    .io_ins_246(rport_io_ins_246),
    .io_ins_247(rport_io_ins_247),
    .io_ins_248(rport_io_ins_248),
    .io_ins_249(rport_io_ins_249),
    .io_ins_250(rport_io_ins_250),
    .io_ins_251(rport_io_ins_251),
    .io_ins_252(rport_io_ins_252),
    .io_ins_253(rport_io_ins_253),
    .io_ins_254(rport_io_ins_254),
    .io_ins_255(rport_io_ins_255),
    .io_ins_256(rport_io_ins_256),
    .io_ins_257(rport_io_ins_257),
    .io_ins_258(rport_io_ins_258),
    .io_ins_259(rport_io_ins_259),
    .io_ins_260(rport_io_ins_260),
    .io_ins_261(rport_io_ins_261),
    .io_ins_262(rport_io_ins_262),
    .io_ins_263(rport_io_ins_263),
    .io_ins_264(rport_io_ins_264),
    .io_ins_265(rport_io_ins_265),
    .io_ins_266(rport_io_ins_266),
    .io_ins_267(rport_io_ins_267),
    .io_ins_268(rport_io_ins_268),
    .io_ins_269(rport_io_ins_269),
    .io_ins_270(rport_io_ins_270),
    .io_ins_271(rport_io_ins_271),
    .io_ins_272(rport_io_ins_272),
    .io_ins_273(rport_io_ins_273),
    .io_ins_274(rport_io_ins_274),
    .io_ins_275(rport_io_ins_275),
    .io_ins_276(rport_io_ins_276),
    .io_ins_277(rport_io_ins_277),
    .io_ins_278(rport_io_ins_278),
    .io_ins_279(rport_io_ins_279),
    .io_ins_280(rport_io_ins_280),
    .io_ins_281(rport_io_ins_281),
    .io_ins_282(rport_io_ins_282),
    .io_ins_283(rport_io_ins_283),
    .io_ins_284(rport_io_ins_284),
    .io_ins_285(rport_io_ins_285),
    .io_ins_286(rport_io_ins_286),
    .io_ins_287(rport_io_ins_287),
    .io_ins_288(rport_io_ins_288),
    .io_ins_289(rport_io_ins_289),
    .io_ins_290(rport_io_ins_290),
    .io_ins_291(rport_io_ins_291),
    .io_ins_292(rport_io_ins_292),
    .io_ins_293(rport_io_ins_293),
    .io_ins_294(rport_io_ins_294),
    .io_ins_295(rport_io_ins_295),
    .io_ins_296(rport_io_ins_296),
    .io_ins_297(rport_io_ins_297),
    .io_ins_298(rport_io_ins_298),
    .io_ins_299(rport_io_ins_299),
    .io_ins_300(rport_io_ins_300),
    .io_ins_301(rport_io_ins_301),
    .io_ins_302(rport_io_ins_302),
    .io_ins_303(rport_io_ins_303),
    .io_ins_304(rport_io_ins_304),
    .io_ins_305(rport_io_ins_305),
    .io_ins_306(rport_io_ins_306),
    .io_ins_307(rport_io_ins_307),
    .io_ins_308(rport_io_ins_308),
    .io_ins_309(rport_io_ins_309),
    .io_ins_310(rport_io_ins_310),
    .io_ins_311(rport_io_ins_311),
    .io_ins_312(rport_io_ins_312),
    .io_ins_313(rport_io_ins_313),
    .io_ins_314(rport_io_ins_314),
    .io_ins_315(rport_io_ins_315),
    .io_ins_316(rport_io_ins_316),
    .io_ins_317(rport_io_ins_317),
    .io_ins_318(rport_io_ins_318),
    .io_ins_319(rport_io_ins_319),
    .io_ins_320(rport_io_ins_320),
    .io_ins_321(rport_io_ins_321),
    .io_ins_322(rport_io_ins_322),
    .io_ins_323(rport_io_ins_323),
    .io_ins_324(rport_io_ins_324),
    .io_ins_325(rport_io_ins_325),
    .io_ins_326(rport_io_ins_326),
    .io_ins_327(rport_io_ins_327),
    .io_ins_328(rport_io_ins_328),
    .io_ins_329(rport_io_ins_329),
    .io_ins_330(rport_io_ins_330),
    .io_ins_331(rport_io_ins_331),
    .io_ins_332(rport_io_ins_332),
    .io_ins_333(rport_io_ins_333),
    .io_ins_334(rport_io_ins_334),
    .io_ins_335(rport_io_ins_335),
    .io_ins_336(rport_io_ins_336),
    .io_ins_337(rport_io_ins_337),
    .io_ins_338(rport_io_ins_338),
    .io_ins_339(rport_io_ins_339),
    .io_ins_340(rport_io_ins_340),
    .io_ins_341(rport_io_ins_341),
    .io_ins_342(rport_io_ins_342),
    .io_ins_343(rport_io_ins_343),
    .io_ins_344(rport_io_ins_344),
    .io_ins_345(rport_io_ins_345),
    .io_ins_346(rport_io_ins_346),
    .io_ins_347(rport_io_ins_347),
    .io_ins_348(rport_io_ins_348),
    .io_ins_349(rport_io_ins_349),
    .io_ins_350(rport_io_ins_350),
    .io_ins_351(rport_io_ins_351),
    .io_ins_352(rport_io_ins_352),
    .io_ins_353(rport_io_ins_353),
    .io_ins_354(rport_io_ins_354),
    .io_ins_355(rport_io_ins_355),
    .io_ins_356(rport_io_ins_356),
    .io_ins_357(rport_io_ins_357),
    .io_ins_358(rport_io_ins_358),
    .io_ins_359(rport_io_ins_359),
    .io_ins_360(rport_io_ins_360),
    .io_ins_361(rport_io_ins_361),
    .io_ins_362(rport_io_ins_362),
    .io_ins_363(rport_io_ins_363),
    .io_ins_364(rport_io_ins_364),
    .io_ins_365(rport_io_ins_365),
    .io_ins_366(rport_io_ins_366),
    .io_ins_367(rport_io_ins_367),
    .io_ins_368(rport_io_ins_368),
    .io_ins_369(rport_io_ins_369),
    .io_ins_370(rport_io_ins_370),
    .io_ins_371(rport_io_ins_371),
    .io_ins_372(rport_io_ins_372),
    .io_ins_373(rport_io_ins_373),
    .io_ins_374(rport_io_ins_374),
    .io_ins_375(rport_io_ins_375),
    .io_ins_376(rport_io_ins_376),
    .io_ins_377(rport_io_ins_377),
    .io_ins_378(rport_io_ins_378),
    .io_ins_379(rport_io_ins_379),
    .io_ins_380(rport_io_ins_380),
    .io_ins_381(rport_io_ins_381),
    .io_ins_382(rport_io_ins_382),
    .io_ins_383(rport_io_ins_383),
    .io_ins_384(rport_io_ins_384),
    .io_ins_385(rport_io_ins_385),
    .io_ins_386(rport_io_ins_386),
    .io_ins_387(rport_io_ins_387),
    .io_ins_388(rport_io_ins_388),
    .io_ins_389(rport_io_ins_389),
    .io_ins_390(rport_io_ins_390),
    .io_ins_391(rport_io_ins_391),
    .io_ins_392(rport_io_ins_392),
    .io_ins_393(rport_io_ins_393),
    .io_ins_394(rport_io_ins_394),
    .io_ins_395(rport_io_ins_395),
    .io_ins_396(rport_io_ins_396),
    .io_ins_397(rport_io_ins_397),
    .io_ins_398(rport_io_ins_398),
    .io_ins_399(rport_io_ins_399),
    .io_ins_400(rport_io_ins_400),
    .io_ins_401(rport_io_ins_401),
    .io_ins_402(rport_io_ins_402),
    .io_ins_403(rport_io_ins_403),
    .io_ins_404(rport_io_ins_404),
    .io_ins_405(rport_io_ins_405),
    .io_ins_406(rport_io_ins_406),
    .io_ins_407(rport_io_ins_407),
    .io_ins_408(rport_io_ins_408),
    .io_ins_409(rport_io_ins_409),
    .io_ins_410(rport_io_ins_410),
    .io_ins_411(rport_io_ins_411),
    .io_ins_412(rport_io_ins_412),
    .io_ins_413(rport_io_ins_413),
    .io_ins_414(rport_io_ins_414),
    .io_ins_415(rport_io_ins_415),
    .io_ins_416(rport_io_ins_416),
    .io_ins_417(rport_io_ins_417),
    .io_ins_418(rport_io_ins_418),
    .io_ins_419(rport_io_ins_419),
    .io_ins_420(rport_io_ins_420),
    .io_ins_421(rport_io_ins_421),
    .io_ins_422(rport_io_ins_422),
    .io_ins_423(rport_io_ins_423),
    .io_ins_424(rport_io_ins_424),
    .io_ins_425(rport_io_ins_425),
    .io_ins_426(rport_io_ins_426),
    .io_ins_427(rport_io_ins_427),
    .io_ins_428(rport_io_ins_428),
    .io_ins_429(rport_io_ins_429),
    .io_ins_430(rport_io_ins_430),
    .io_ins_431(rport_io_ins_431),
    .io_ins_432(rport_io_ins_432),
    .io_ins_433(rport_io_ins_433),
    .io_ins_434(rport_io_ins_434),
    .io_ins_435(rport_io_ins_435),
    .io_ins_436(rport_io_ins_436),
    .io_ins_437(rport_io_ins_437),
    .io_ins_438(rport_io_ins_438),
    .io_ins_439(rport_io_ins_439),
    .io_ins_440(rport_io_ins_440),
    .io_ins_441(rport_io_ins_441),
    .io_ins_442(rport_io_ins_442),
    .io_ins_443(rport_io_ins_443),
    .io_ins_444(rport_io_ins_444),
    .io_ins_445(rport_io_ins_445),
    .io_ins_446(rport_io_ins_446),
    .io_ins_447(rport_io_ins_447),
    .io_ins_448(rport_io_ins_448),
    .io_ins_449(rport_io_ins_449),
    .io_ins_450(rport_io_ins_450),
    .io_ins_451(rport_io_ins_451),
    .io_ins_452(rport_io_ins_452),
    .io_ins_453(rport_io_ins_453),
    .io_ins_454(rport_io_ins_454),
    .io_ins_455(rport_io_ins_455),
    .io_ins_456(rport_io_ins_456),
    .io_ins_457(rport_io_ins_457),
    .io_ins_458(rport_io_ins_458),
    .io_ins_459(rport_io_ins_459),
    .io_ins_460(rport_io_ins_460),
    .io_ins_461(rport_io_ins_461),
    .io_ins_462(rport_io_ins_462),
    .io_ins_463(rport_io_ins_463),
    .io_ins_464(rport_io_ins_464),
    .io_ins_465(rport_io_ins_465),
    .io_ins_466(rport_io_ins_466),
    .io_ins_467(rport_io_ins_467),
    .io_ins_468(rport_io_ins_468),
    .io_ins_469(rport_io_ins_469),
    .io_ins_470(rport_io_ins_470),
    .io_ins_471(rport_io_ins_471),
    .io_ins_472(rport_io_ins_472),
    .io_ins_473(rport_io_ins_473),
    .io_ins_474(rport_io_ins_474),
    .io_ins_475(rport_io_ins_475),
    .io_ins_476(rport_io_ins_476),
    .io_ins_477(rport_io_ins_477),
    .io_ins_478(rport_io_ins_478),
    .io_ins_479(rport_io_ins_479),
    .io_ins_480(rport_io_ins_480),
    .io_ins_481(rport_io_ins_481),
    .io_ins_482(rport_io_ins_482),
    .io_ins_483(rport_io_ins_483),
    .io_ins_484(rport_io_ins_484),
    .io_ins_485(rport_io_ins_485),
    .io_ins_486(rport_io_ins_486),
    .io_ins_487(rport_io_ins_487),
    .io_ins_488(rport_io_ins_488),
    .io_ins_489(rport_io_ins_489),
    .io_ins_490(rport_io_ins_490),
    .io_ins_491(rport_io_ins_491),
    .io_ins_492(rport_io_ins_492),
    .io_ins_493(rport_io_ins_493),
    .io_ins_494(rport_io_ins_494),
    .io_ins_495(rport_io_ins_495),
    .io_ins_496(rport_io_ins_496),
    .io_ins_497(rport_io_ins_497),
    .io_ins_498(rport_io_ins_498),
    .io_ins_499(rport_io_ins_499),
    .io_ins_500(rport_io_ins_500),
    .io_ins_501(rport_io_ins_501),
    .io_ins_502(rport_io_ins_502),
    .io_ins_503(rport_io_ins_503),
    .io_ins_504(rport_io_ins_504),
    .io_ins_505(rport_io_ins_505),
    .io_sel(rport_io_sel),
    .io_out(rport_io_out)
  );
  assign _T_1544 = io_waddr == 32'h0;
  assign _T_1545 = io_wen & _T_1544;
  assign _T_1550 = io_waddr == 32'h1;
  assign _T_1551 = io_wen & _T_1550;
  assign _T_1555 = _T_1551 ? _T_1551 : io_argOuts_0_valid;
  assign _T_1559 = _T_1551 ? io_wdata : io_argOuts_0_bits;
  assign _T_1564 = io_waddr == 32'h2;
  assign _T_1565 = io_wen & _T_1564;
  assign _T_1570 = io_waddr == 32'h3;
  assign _T_1571 = io_wen & _T_1570;
  assign _T_1576 = io_waddr == 32'h4;
  assign _T_1577 = io_wen & _T_1576;
  assign _T_1582 = io_waddr == 32'h5;
  assign _T_1583 = io_wen & _T_1582;
  assign _T_1584 = io_argOuts_1_valid | _T_1583;
  assign _T_1585 = io_argOuts_1_valid ? io_argOuts_1_bits : io_wdata;
  assign _T_5611 = io_raddr & 32'hfffeffff;
  assign _T_5612 = io_raddr[16];
  assign _T_5613 = rport_io_out[63:32];
  assign _T_5614 = rport_io_out[31:0];
  assign _T_5615 = _T_5612 ? _T_5613 : _T_5614;
  assign io_rdata = {{32'd0}, _T_5615};
  assign io_argIns_0 = _T_5618_0;
  assign io_argIns_1 = _T_5618_1;
  assign io_argIns_2 = _T_5618_2;
  assign io_argIns_3 = _T_5618_3;
  assign io_argIns_4 = _T_5618_4;
  assign regs_0_io_in = io_wdata;
  assign regs_0_io_init = 64'h0;
  assign regs_0_io_reset = reset;
  assign regs_0_io_enable = _T_1545;
  assign regs_0_clock = clock;
  assign regs_0_reset = reset;
  assign regs_1_io_in = _T_1559;
  assign regs_1_io_init = 64'h0;
  assign regs_1_io_reset = reset;
  assign regs_1_io_enable = _T_1555;
  assign regs_1_clock = clock;
  assign regs_1_reset = reset;
  assign regs_2_io_in = io_wdata;
  assign regs_2_io_init = 64'h0;
  assign regs_2_io_reset = reset;
  assign regs_2_io_enable = _T_1565;
  assign regs_2_clock = clock;
  assign regs_2_reset = reset;
  assign regs_3_io_in = io_wdata;
  assign regs_3_io_init = 64'h0;
  assign regs_3_io_reset = reset;
  assign regs_3_io_enable = _T_1571;
  assign regs_3_clock = clock;
  assign regs_3_reset = reset;
  assign regs_4_io_in = io_wdata;
  assign regs_4_io_init = 64'h0;
  assign regs_4_io_reset = reset;
  assign regs_4_io_enable = _T_1577;
  assign regs_4_clock = clock;
  assign regs_4_reset = reset;
  assign regs_5_io_in = _T_1585;
  assign regs_5_io_init = 64'h0;
  assign regs_5_io_reset = reset;
  assign regs_5_io_enable = _T_1584;
  assign regs_5_clock = clock;
  assign regs_5_reset = io_reset;
  assign regs_6_io_in = io_argOuts_2_bits;
  assign regs_6_io_init = 64'h0;
  assign regs_6_io_reset = reset;
  assign regs_6_io_enable = 1'h1;
  assign regs_6_clock = clock;
  assign regs_6_reset = io_reset;
  assign regs_7_io_in = io_argOuts_3_bits;
  assign regs_7_io_init = 64'h0;
  assign regs_7_io_reset = reset;
  assign regs_7_io_enable = 1'h1;
  assign regs_7_clock = clock;
  assign regs_7_reset = io_reset;
  assign regs_8_io_in = io_argOuts_4_bits;
  assign regs_8_io_init = 64'h0;
  assign regs_8_io_reset = reset;
  assign regs_8_io_enable = 1'h1;
  assign regs_8_clock = clock;
  assign regs_8_reset = io_reset;
  assign regs_9_io_in = io_argOuts_5_bits;
  assign regs_9_io_init = 64'h0;
  assign regs_9_io_reset = reset;
  assign regs_9_io_enable = 1'h1;
  assign regs_9_clock = clock;
  assign regs_9_reset = io_reset;
  assign regs_10_io_in = io_argOuts_6_bits;
  assign regs_10_io_init = 64'h0;
  assign regs_10_io_reset = reset;
  assign regs_10_io_enable = 1'h1;
  assign regs_10_clock = clock;
  assign regs_10_reset = io_reset;
  assign regs_11_io_in = io_argOuts_7_bits;
  assign regs_11_io_init = 64'h0;
  assign regs_11_io_reset = reset;
  assign regs_11_io_enable = 1'h1;
  assign regs_11_clock = clock;
  assign regs_11_reset = io_reset;
  assign regs_12_io_in = io_argOuts_8_bits;
  assign regs_12_io_init = 64'h0;
  assign regs_12_io_reset = reset;
  assign regs_12_io_enable = 1'h1;
  assign regs_12_clock = clock;
  assign regs_12_reset = io_reset;
  assign regs_13_io_in = io_argOuts_9_bits;
  assign regs_13_io_init = 64'h0;
  assign regs_13_io_reset = reset;
  assign regs_13_io_enable = 1'h1;
  assign regs_13_clock = clock;
  assign regs_13_reset = io_reset;
  assign regs_14_io_in = io_argOuts_10_bits;
  assign regs_14_io_init = 64'h0;
  assign regs_14_io_reset = reset;
  assign regs_14_io_enable = 1'h1;
  assign regs_14_clock = clock;
  assign regs_14_reset = io_reset;
  assign regs_15_io_in = io_argOuts_11_bits;
  assign regs_15_io_init = 64'h0;
  assign regs_15_io_reset = reset;
  assign regs_15_io_enable = 1'h1;
  assign regs_15_clock = clock;
  assign regs_15_reset = io_reset;
  assign regs_16_io_in = io_argOuts_12_bits;
  assign regs_16_io_init = 64'h0;
  assign regs_16_io_reset = reset;
  assign regs_16_io_enable = 1'h1;
  assign regs_16_clock = clock;
  assign regs_16_reset = io_reset;
  assign regs_17_io_in = io_argOuts_13_bits;
  assign regs_17_io_init = 64'h0;
  assign regs_17_io_reset = reset;
  assign regs_17_io_enable = 1'h1;
  assign regs_17_clock = clock;
  assign regs_17_reset = io_reset;
  assign regs_18_io_in = io_argOuts_14_bits;
  assign regs_18_io_init = 64'h0;
  assign regs_18_io_reset = reset;
  assign regs_18_io_enable = 1'h1;
  assign regs_18_clock = clock;
  assign regs_18_reset = io_reset;
  assign regs_19_io_in = io_argOuts_15_bits;
  assign regs_19_io_init = 64'h0;
  assign regs_19_io_reset = reset;
  assign regs_19_io_enable = 1'h1;
  assign regs_19_clock = clock;
  assign regs_19_reset = io_reset;
  assign regs_20_io_in = io_argOuts_16_bits;
  assign regs_20_io_init = 64'h0;
  assign regs_20_io_reset = reset;
  assign regs_20_io_enable = 1'h1;
  assign regs_20_clock = clock;
  assign regs_20_reset = io_reset;
  assign regs_21_io_in = io_argOuts_17_bits;
  assign regs_21_io_init = 64'h0;
  assign regs_21_io_reset = reset;
  assign regs_21_io_enable = 1'h1;
  assign regs_21_clock = clock;
  assign regs_21_reset = io_reset;
  assign regs_22_io_in = io_argOuts_18_bits;
  assign regs_22_io_init = 64'h0;
  assign regs_22_io_reset = reset;
  assign regs_22_io_enable = 1'h1;
  assign regs_22_clock = clock;
  assign regs_22_reset = io_reset;
  assign regs_23_io_in = io_argOuts_19_bits;
  assign regs_23_io_init = 64'h0;
  assign regs_23_io_reset = reset;
  assign regs_23_io_enable = 1'h1;
  assign regs_23_clock = clock;
  assign regs_23_reset = io_reset;
  assign regs_24_io_in = io_argOuts_20_bits;
  assign regs_24_io_init = 64'h0;
  assign regs_24_io_reset = reset;
  assign regs_24_io_enable = 1'h1;
  assign regs_24_clock = clock;
  assign regs_24_reset = io_reset;
  assign regs_25_io_in = io_argOuts_21_bits;
  assign regs_25_io_init = 64'h0;
  assign regs_25_io_reset = reset;
  assign regs_25_io_enable = 1'h1;
  assign regs_25_clock = clock;
  assign regs_25_reset = io_reset;
  assign regs_26_io_in = io_argOuts_22_bits;
  assign regs_26_io_init = 64'h0;
  assign regs_26_io_reset = reset;
  assign regs_26_io_enable = 1'h1;
  assign regs_26_clock = clock;
  assign regs_26_reset = io_reset;
  assign regs_27_io_in = io_argOuts_23_bits;
  assign regs_27_io_init = 64'h0;
  assign regs_27_io_reset = reset;
  assign regs_27_io_enable = 1'h1;
  assign regs_27_clock = clock;
  assign regs_27_reset = io_reset;
  assign regs_28_io_in = io_argOuts_24_bits;
  assign regs_28_io_init = 64'h0;
  assign regs_28_io_reset = reset;
  assign regs_28_io_enable = 1'h1;
  assign regs_28_clock = clock;
  assign regs_28_reset = io_reset;
  assign regs_29_io_in = io_argOuts_25_bits;
  assign regs_29_io_init = 64'h0;
  assign regs_29_io_reset = reset;
  assign regs_29_io_enable = 1'h1;
  assign regs_29_clock = clock;
  assign regs_29_reset = io_reset;
  assign regs_30_io_in = io_argOuts_26_bits;
  assign regs_30_io_init = 64'h0;
  assign regs_30_io_reset = reset;
  assign regs_30_io_enable = 1'h1;
  assign regs_30_clock = clock;
  assign regs_30_reset = io_reset;
  assign regs_31_io_in = io_argOuts_27_bits;
  assign regs_31_io_init = 64'h0;
  assign regs_31_io_reset = reset;
  assign regs_31_io_enable = 1'h1;
  assign regs_31_clock = clock;
  assign regs_31_reset = io_reset;
  assign regs_32_io_in = io_argOuts_28_bits;
  assign regs_32_io_init = 64'h0;
  assign regs_32_io_reset = reset;
  assign regs_32_io_enable = 1'h1;
  assign regs_32_clock = clock;
  assign regs_32_reset = io_reset;
  assign regs_33_io_in = io_argOuts_29_bits;
  assign regs_33_io_init = 64'h0;
  assign regs_33_io_reset = reset;
  assign regs_33_io_enable = 1'h1;
  assign regs_33_clock = clock;
  assign regs_33_reset = io_reset;
  assign regs_34_io_in = io_argOuts_30_bits;
  assign regs_34_io_init = 64'h0;
  assign regs_34_io_reset = reset;
  assign regs_34_io_enable = 1'h1;
  assign regs_34_clock = clock;
  assign regs_34_reset = io_reset;
  assign regs_35_io_in = io_argOuts_31_bits;
  assign regs_35_io_init = 64'h0;
  assign regs_35_io_reset = reset;
  assign regs_35_io_enable = 1'h1;
  assign regs_35_clock = clock;
  assign regs_35_reset = io_reset;
  assign regs_36_io_in = io_argOuts_32_bits;
  assign regs_36_io_init = 64'h0;
  assign regs_36_io_reset = reset;
  assign regs_36_io_enable = 1'h1;
  assign regs_36_clock = clock;
  assign regs_36_reset = io_reset;
  assign regs_37_io_in = io_argOuts_33_bits;
  assign regs_37_io_init = 64'h0;
  assign regs_37_io_reset = reset;
  assign regs_37_io_enable = 1'h1;
  assign regs_37_clock = clock;
  assign regs_37_reset = io_reset;
  assign regs_38_io_in = io_argOuts_34_bits;
  assign regs_38_io_init = 64'h0;
  assign regs_38_io_reset = reset;
  assign regs_38_io_enable = 1'h1;
  assign regs_38_clock = clock;
  assign regs_38_reset = io_reset;
  assign regs_39_io_in = io_argOuts_35_bits;
  assign regs_39_io_init = 64'h0;
  assign regs_39_io_reset = reset;
  assign regs_39_io_enable = 1'h1;
  assign regs_39_clock = clock;
  assign regs_39_reset = io_reset;
  assign regs_40_io_in = io_argOuts_36_bits;
  assign regs_40_io_init = 64'h0;
  assign regs_40_io_reset = reset;
  assign regs_40_io_enable = 1'h1;
  assign regs_40_clock = clock;
  assign regs_40_reset = io_reset;
  assign regs_41_io_in = io_argOuts_37_bits;
  assign regs_41_io_init = 64'h0;
  assign regs_41_io_reset = reset;
  assign regs_41_io_enable = 1'h1;
  assign regs_41_clock = clock;
  assign regs_41_reset = io_reset;
  assign regs_42_io_in = io_argOuts_38_bits;
  assign regs_42_io_init = 64'h0;
  assign regs_42_io_reset = reset;
  assign regs_42_io_enable = 1'h1;
  assign regs_42_clock = clock;
  assign regs_42_reset = io_reset;
  assign regs_43_io_in = io_argOuts_39_bits;
  assign regs_43_io_init = 64'h0;
  assign regs_43_io_reset = reset;
  assign regs_43_io_enable = 1'h1;
  assign regs_43_clock = clock;
  assign regs_43_reset = io_reset;
  assign regs_44_io_in = io_argOuts_40_bits;
  assign regs_44_io_init = 64'h0;
  assign regs_44_io_reset = reset;
  assign regs_44_io_enable = 1'h1;
  assign regs_44_clock = clock;
  assign regs_44_reset = io_reset;
  assign regs_45_io_in = io_argOuts_41_bits;
  assign regs_45_io_init = 64'h0;
  assign regs_45_io_reset = reset;
  assign regs_45_io_enable = 1'h1;
  assign regs_45_clock = clock;
  assign regs_45_reset = io_reset;
  assign regs_46_io_in = io_argOuts_42_bits;
  assign regs_46_io_init = 64'h0;
  assign regs_46_io_reset = reset;
  assign regs_46_io_enable = 1'h1;
  assign regs_46_clock = clock;
  assign regs_46_reset = io_reset;
  assign regs_47_io_in = io_argOuts_43_bits;
  assign regs_47_io_init = 64'h0;
  assign regs_47_io_reset = reset;
  assign regs_47_io_enable = 1'h1;
  assign regs_47_clock = clock;
  assign regs_47_reset = io_reset;
  assign regs_48_io_in = io_argOuts_44_bits;
  assign regs_48_io_init = 64'h0;
  assign regs_48_io_reset = reset;
  assign regs_48_io_enable = 1'h1;
  assign regs_48_clock = clock;
  assign regs_48_reset = io_reset;
  assign regs_49_io_in = io_argOuts_45_bits;
  assign regs_49_io_init = 64'h0;
  assign regs_49_io_reset = reset;
  assign regs_49_io_enable = 1'h1;
  assign regs_49_clock = clock;
  assign regs_49_reset = io_reset;
  assign regs_50_io_in = io_argOuts_46_bits;
  assign regs_50_io_init = 64'h0;
  assign regs_50_io_reset = reset;
  assign regs_50_io_enable = 1'h1;
  assign regs_50_clock = clock;
  assign regs_50_reset = io_reset;
  assign regs_51_io_in = io_argOuts_47_bits;
  assign regs_51_io_init = 64'h0;
  assign regs_51_io_reset = reset;
  assign regs_51_io_enable = 1'h1;
  assign regs_51_clock = clock;
  assign regs_51_reset = io_reset;
  assign regs_52_io_in = io_argOuts_48_bits;
  assign regs_52_io_init = 64'h0;
  assign regs_52_io_reset = reset;
  assign regs_52_io_enable = 1'h1;
  assign regs_52_clock = clock;
  assign regs_52_reset = io_reset;
  assign regs_53_io_in = io_argOuts_49_bits;
  assign regs_53_io_init = 64'h0;
  assign regs_53_io_reset = reset;
  assign regs_53_io_enable = 1'h1;
  assign regs_53_clock = clock;
  assign regs_53_reset = io_reset;
  assign regs_54_io_in = io_argOuts_50_bits;
  assign regs_54_io_init = 64'h0;
  assign regs_54_io_reset = reset;
  assign regs_54_io_enable = 1'h1;
  assign regs_54_clock = clock;
  assign regs_54_reset = io_reset;
  assign regs_55_io_in = io_argOuts_51_bits;
  assign regs_55_io_init = 64'h0;
  assign regs_55_io_reset = reset;
  assign regs_55_io_enable = 1'h1;
  assign regs_55_clock = clock;
  assign regs_55_reset = io_reset;
  assign regs_56_io_in = io_argOuts_52_bits;
  assign regs_56_io_init = 64'h0;
  assign regs_56_io_reset = reset;
  assign regs_56_io_enable = 1'h1;
  assign regs_56_clock = clock;
  assign regs_56_reset = io_reset;
  assign regs_57_io_in = io_argOuts_53_bits;
  assign regs_57_io_init = 64'h0;
  assign regs_57_io_reset = reset;
  assign regs_57_io_enable = 1'h1;
  assign regs_57_clock = clock;
  assign regs_57_reset = io_reset;
  assign regs_58_io_in = io_argOuts_54_bits;
  assign regs_58_io_init = 64'h0;
  assign regs_58_io_reset = reset;
  assign regs_58_io_enable = 1'h1;
  assign regs_58_clock = clock;
  assign regs_58_reset = io_reset;
  assign regs_59_io_in = io_argOuts_55_bits;
  assign regs_59_io_init = 64'h0;
  assign regs_59_io_reset = reset;
  assign regs_59_io_enable = 1'h1;
  assign regs_59_clock = clock;
  assign regs_59_reset = io_reset;
  assign regs_60_io_in = io_argOuts_56_bits;
  assign regs_60_io_init = 64'h0;
  assign regs_60_io_reset = reset;
  assign regs_60_io_enable = 1'h1;
  assign regs_60_clock = clock;
  assign regs_60_reset = io_reset;
  assign regs_61_io_in = io_argOuts_57_bits;
  assign regs_61_io_init = 64'h0;
  assign regs_61_io_reset = reset;
  assign regs_61_io_enable = 1'h1;
  assign regs_61_clock = clock;
  assign regs_61_reset = io_reset;
  assign regs_62_io_in = io_argOuts_58_bits;
  assign regs_62_io_init = 64'h0;
  assign regs_62_io_reset = reset;
  assign regs_62_io_enable = 1'h1;
  assign regs_62_clock = clock;
  assign regs_62_reset = io_reset;
  assign regs_63_io_in = io_argOuts_59_bits;
  assign regs_63_io_init = 64'h0;
  assign regs_63_io_reset = reset;
  assign regs_63_io_enable = 1'h1;
  assign regs_63_clock = clock;
  assign regs_63_reset = io_reset;
  assign regs_64_io_in = io_argOuts_60_bits;
  assign regs_64_io_init = 64'h0;
  assign regs_64_io_reset = reset;
  assign regs_64_io_enable = 1'h1;
  assign regs_64_clock = clock;
  assign regs_64_reset = io_reset;
  assign regs_65_io_in = io_argOuts_61_bits;
  assign regs_65_io_init = 64'h0;
  assign regs_65_io_reset = reset;
  assign regs_65_io_enable = 1'h1;
  assign regs_65_clock = clock;
  assign regs_65_reset = io_reset;
  assign regs_66_io_in = io_argOuts_62_bits;
  assign regs_66_io_init = 64'h0;
  assign regs_66_io_reset = reset;
  assign regs_66_io_enable = 1'h1;
  assign regs_66_clock = clock;
  assign regs_66_reset = io_reset;
  assign regs_67_io_in = io_argOuts_63_bits;
  assign regs_67_io_init = 64'h0;
  assign regs_67_io_reset = reset;
  assign regs_67_io_enable = 1'h1;
  assign regs_67_clock = clock;
  assign regs_67_reset = io_reset;
  assign regs_68_io_in = io_argOuts_64_bits;
  assign regs_68_io_init = 64'h0;
  assign regs_68_io_reset = reset;
  assign regs_68_io_enable = 1'h1;
  assign regs_68_clock = clock;
  assign regs_68_reset = io_reset;
  assign regs_69_io_in = io_argOuts_65_bits;
  assign regs_69_io_init = 64'h0;
  assign regs_69_io_reset = reset;
  assign regs_69_io_enable = 1'h1;
  assign regs_69_clock = clock;
  assign regs_69_reset = io_reset;
  assign regs_70_io_in = io_argOuts_66_bits;
  assign regs_70_io_init = 64'h0;
  assign regs_70_io_reset = reset;
  assign regs_70_io_enable = 1'h1;
  assign regs_70_clock = clock;
  assign regs_70_reset = io_reset;
  assign regs_71_io_in = io_argOuts_67_bits;
  assign regs_71_io_init = 64'h0;
  assign regs_71_io_reset = reset;
  assign regs_71_io_enable = 1'h1;
  assign regs_71_clock = clock;
  assign regs_71_reset = io_reset;
  assign regs_72_io_in = io_argOuts_68_bits;
  assign regs_72_io_init = 64'h0;
  assign regs_72_io_reset = reset;
  assign regs_72_io_enable = 1'h1;
  assign regs_72_clock = clock;
  assign regs_72_reset = io_reset;
  assign regs_73_io_in = io_argOuts_69_bits;
  assign regs_73_io_init = 64'h0;
  assign regs_73_io_reset = reset;
  assign regs_73_io_enable = 1'h1;
  assign regs_73_clock = clock;
  assign regs_73_reset = io_reset;
  assign regs_74_io_in = io_argOuts_70_bits;
  assign regs_74_io_init = 64'h0;
  assign regs_74_io_reset = reset;
  assign regs_74_io_enable = 1'h1;
  assign regs_74_clock = clock;
  assign regs_74_reset = io_reset;
  assign regs_75_io_in = io_argOuts_71_bits;
  assign regs_75_io_init = 64'h0;
  assign regs_75_io_reset = reset;
  assign regs_75_io_enable = 1'h1;
  assign regs_75_clock = clock;
  assign regs_75_reset = io_reset;
  assign regs_76_io_in = io_argOuts_72_bits;
  assign regs_76_io_init = 64'h0;
  assign regs_76_io_reset = reset;
  assign regs_76_io_enable = 1'h1;
  assign regs_76_clock = clock;
  assign regs_76_reset = io_reset;
  assign regs_77_io_in = io_argOuts_73_bits;
  assign regs_77_io_init = 64'h0;
  assign regs_77_io_reset = reset;
  assign regs_77_io_enable = 1'h1;
  assign regs_77_clock = clock;
  assign regs_77_reset = io_reset;
  assign regs_78_io_in = io_argOuts_74_bits;
  assign regs_78_io_init = 64'h0;
  assign regs_78_io_reset = reset;
  assign regs_78_io_enable = 1'h1;
  assign regs_78_clock = clock;
  assign regs_78_reset = io_reset;
  assign regs_79_io_in = io_argOuts_75_bits;
  assign regs_79_io_init = 64'h0;
  assign regs_79_io_reset = reset;
  assign regs_79_io_enable = 1'h1;
  assign regs_79_clock = clock;
  assign regs_79_reset = io_reset;
  assign regs_80_io_in = io_argOuts_76_bits;
  assign regs_80_io_init = 64'h0;
  assign regs_80_io_reset = reset;
  assign regs_80_io_enable = 1'h1;
  assign regs_80_clock = clock;
  assign regs_80_reset = io_reset;
  assign regs_81_io_in = io_argOuts_77_bits;
  assign regs_81_io_init = 64'h0;
  assign regs_81_io_reset = reset;
  assign regs_81_io_enable = 1'h1;
  assign regs_81_clock = clock;
  assign regs_81_reset = io_reset;
  assign regs_82_io_in = io_argOuts_78_bits;
  assign regs_82_io_init = 64'h0;
  assign regs_82_io_reset = reset;
  assign regs_82_io_enable = 1'h1;
  assign regs_82_clock = clock;
  assign regs_82_reset = io_reset;
  assign regs_83_io_in = io_argOuts_79_bits;
  assign regs_83_io_init = 64'h0;
  assign regs_83_io_reset = reset;
  assign regs_83_io_enable = 1'h1;
  assign regs_83_clock = clock;
  assign regs_83_reset = io_reset;
  assign regs_84_io_in = io_argOuts_80_bits;
  assign regs_84_io_init = 64'h0;
  assign regs_84_io_reset = reset;
  assign regs_84_io_enable = 1'h1;
  assign regs_84_clock = clock;
  assign regs_84_reset = io_reset;
  assign regs_85_io_in = io_argOuts_81_bits;
  assign regs_85_io_init = 64'h0;
  assign regs_85_io_reset = reset;
  assign regs_85_io_enable = 1'h1;
  assign regs_85_clock = clock;
  assign regs_85_reset = io_reset;
  assign regs_86_io_in = io_argOuts_82_bits;
  assign regs_86_io_init = 64'h0;
  assign regs_86_io_reset = reset;
  assign regs_86_io_enable = 1'h1;
  assign regs_86_clock = clock;
  assign regs_86_reset = io_reset;
  assign regs_87_io_in = io_argOuts_83_bits;
  assign regs_87_io_init = 64'h0;
  assign regs_87_io_reset = reset;
  assign regs_87_io_enable = 1'h1;
  assign regs_87_clock = clock;
  assign regs_87_reset = io_reset;
  assign regs_88_io_in = io_argOuts_84_bits;
  assign regs_88_io_init = 64'h0;
  assign regs_88_io_reset = reset;
  assign regs_88_io_enable = 1'h1;
  assign regs_88_clock = clock;
  assign regs_88_reset = io_reset;
  assign regs_89_io_in = io_argOuts_85_bits;
  assign regs_89_io_init = 64'h0;
  assign regs_89_io_reset = reset;
  assign regs_89_io_enable = 1'h1;
  assign regs_89_clock = clock;
  assign regs_89_reset = io_reset;
  assign regs_90_io_in = io_argOuts_86_bits;
  assign regs_90_io_init = 64'h0;
  assign regs_90_io_reset = reset;
  assign regs_90_io_enable = 1'h1;
  assign regs_90_clock = clock;
  assign regs_90_reset = io_reset;
  assign regs_91_io_in = io_argOuts_87_bits;
  assign regs_91_io_init = 64'h0;
  assign regs_91_io_reset = reset;
  assign regs_91_io_enable = 1'h1;
  assign regs_91_clock = clock;
  assign regs_91_reset = io_reset;
  assign regs_92_io_in = io_argOuts_88_bits;
  assign regs_92_io_init = 64'h0;
  assign regs_92_io_reset = reset;
  assign regs_92_io_enable = 1'h1;
  assign regs_92_clock = clock;
  assign regs_92_reset = io_reset;
  assign regs_93_io_in = io_argOuts_89_bits;
  assign regs_93_io_init = 64'h0;
  assign regs_93_io_reset = reset;
  assign regs_93_io_enable = 1'h1;
  assign regs_93_clock = clock;
  assign regs_93_reset = io_reset;
  assign regs_94_io_in = io_argOuts_90_bits;
  assign regs_94_io_init = 64'h0;
  assign regs_94_io_reset = reset;
  assign regs_94_io_enable = 1'h1;
  assign regs_94_clock = clock;
  assign regs_94_reset = io_reset;
  assign regs_95_io_in = io_argOuts_91_bits;
  assign regs_95_io_init = 64'h0;
  assign regs_95_io_reset = reset;
  assign regs_95_io_enable = 1'h1;
  assign regs_95_clock = clock;
  assign regs_95_reset = io_reset;
  assign regs_96_io_in = io_argOuts_92_bits;
  assign regs_96_io_init = 64'h0;
  assign regs_96_io_reset = reset;
  assign regs_96_io_enable = 1'h1;
  assign regs_96_clock = clock;
  assign regs_96_reset = io_reset;
  assign regs_97_io_in = io_argOuts_93_bits;
  assign regs_97_io_init = 64'h0;
  assign regs_97_io_reset = reset;
  assign regs_97_io_enable = 1'h1;
  assign regs_97_clock = clock;
  assign regs_97_reset = io_reset;
  assign regs_98_io_in = io_argOuts_94_bits;
  assign regs_98_io_init = 64'h0;
  assign regs_98_io_reset = reset;
  assign regs_98_io_enable = 1'h1;
  assign regs_98_clock = clock;
  assign regs_98_reset = io_reset;
  assign regs_99_io_in = io_argOuts_95_bits;
  assign regs_99_io_init = 64'h0;
  assign regs_99_io_reset = reset;
  assign regs_99_io_enable = 1'h1;
  assign regs_99_clock = clock;
  assign regs_99_reset = io_reset;
  assign regs_100_io_in = io_argOuts_96_bits;
  assign regs_100_io_init = 64'h0;
  assign regs_100_io_reset = reset;
  assign regs_100_io_enable = 1'h1;
  assign regs_100_clock = clock;
  assign regs_100_reset = io_reset;
  assign regs_101_io_in = io_argOuts_97_bits;
  assign regs_101_io_init = 64'h0;
  assign regs_101_io_reset = reset;
  assign regs_101_io_enable = 1'h1;
  assign regs_101_clock = clock;
  assign regs_101_reset = io_reset;
  assign regs_102_io_in = io_argOuts_98_bits;
  assign regs_102_io_init = 64'h0;
  assign regs_102_io_reset = reset;
  assign regs_102_io_enable = 1'h1;
  assign regs_102_clock = clock;
  assign regs_102_reset = io_reset;
  assign regs_103_io_in = io_argOuts_99_bits;
  assign regs_103_io_init = 64'h0;
  assign regs_103_io_reset = reset;
  assign regs_103_io_enable = 1'h1;
  assign regs_103_clock = clock;
  assign regs_103_reset = io_reset;
  assign regs_104_io_in = io_argOuts_100_bits;
  assign regs_104_io_init = 64'h0;
  assign regs_104_io_reset = reset;
  assign regs_104_io_enable = 1'h1;
  assign regs_104_clock = clock;
  assign regs_104_reset = io_reset;
  assign regs_105_io_in = io_argOuts_101_bits;
  assign regs_105_io_init = 64'h0;
  assign regs_105_io_reset = reset;
  assign regs_105_io_enable = 1'h1;
  assign regs_105_clock = clock;
  assign regs_105_reset = io_reset;
  assign regs_106_io_in = io_argOuts_102_bits;
  assign regs_106_io_init = 64'h0;
  assign regs_106_io_reset = reset;
  assign regs_106_io_enable = 1'h1;
  assign regs_106_clock = clock;
  assign regs_106_reset = io_reset;
  assign regs_107_io_in = io_argOuts_103_bits;
  assign regs_107_io_init = 64'h0;
  assign regs_107_io_reset = reset;
  assign regs_107_io_enable = 1'h1;
  assign regs_107_clock = clock;
  assign regs_107_reset = io_reset;
  assign regs_108_io_in = io_argOuts_104_bits;
  assign regs_108_io_init = 64'h0;
  assign regs_108_io_reset = reset;
  assign regs_108_io_enable = 1'h1;
  assign regs_108_clock = clock;
  assign regs_108_reset = io_reset;
  assign regs_109_io_in = io_argOuts_105_bits;
  assign regs_109_io_init = 64'h0;
  assign regs_109_io_reset = reset;
  assign regs_109_io_enable = 1'h1;
  assign regs_109_clock = clock;
  assign regs_109_reset = io_reset;
  assign regs_110_io_in = io_argOuts_106_bits;
  assign regs_110_io_init = 64'h0;
  assign regs_110_io_reset = reset;
  assign regs_110_io_enable = 1'h1;
  assign regs_110_clock = clock;
  assign regs_110_reset = io_reset;
  assign regs_111_io_in = io_argOuts_107_bits;
  assign regs_111_io_init = 64'h0;
  assign regs_111_io_reset = reset;
  assign regs_111_io_enable = 1'h1;
  assign regs_111_clock = clock;
  assign regs_111_reset = io_reset;
  assign regs_112_io_in = io_argOuts_108_bits;
  assign regs_112_io_init = 64'h0;
  assign regs_112_io_reset = reset;
  assign regs_112_io_enable = 1'h1;
  assign regs_112_clock = clock;
  assign regs_112_reset = io_reset;
  assign regs_113_io_in = io_argOuts_109_bits;
  assign regs_113_io_init = 64'h0;
  assign regs_113_io_reset = reset;
  assign regs_113_io_enable = 1'h1;
  assign regs_113_clock = clock;
  assign regs_113_reset = io_reset;
  assign regs_114_io_in = 64'h0;
  assign regs_114_io_init = 64'h0;
  assign regs_114_io_reset = reset;
  assign regs_114_io_enable = 1'h1;
  assign regs_114_clock = clock;
  assign regs_114_reset = io_reset;
  assign regs_115_io_in = 64'h0;
  assign regs_115_io_init = 64'h0;
  assign regs_115_io_reset = reset;
  assign regs_115_io_enable = 1'h1;
  assign regs_115_clock = clock;
  assign regs_115_reset = io_reset;
  assign regs_116_io_in = 64'h0;
  assign regs_116_io_init = 64'h0;
  assign regs_116_io_reset = reset;
  assign regs_116_io_enable = 1'h1;
  assign regs_116_clock = clock;
  assign regs_116_reset = io_reset;
  assign regs_117_io_in = 64'h0;
  assign regs_117_io_init = 64'h0;
  assign regs_117_io_reset = reset;
  assign regs_117_io_enable = 1'h1;
  assign regs_117_clock = clock;
  assign regs_117_reset = io_reset;
  assign regs_118_io_in = 64'h0;
  assign regs_118_io_init = 64'h0;
  assign regs_118_io_reset = reset;
  assign regs_118_io_enable = 1'h1;
  assign regs_118_clock = clock;
  assign regs_118_reset = io_reset;
  assign regs_119_io_in = 64'h0;
  assign regs_119_io_init = 64'h0;
  assign regs_119_io_reset = reset;
  assign regs_119_io_enable = 1'h1;
  assign regs_119_clock = clock;
  assign regs_119_reset = io_reset;
  assign regs_120_io_in = 64'h0;
  assign regs_120_io_init = 64'h0;
  assign regs_120_io_reset = reset;
  assign regs_120_io_enable = 1'h1;
  assign regs_120_clock = clock;
  assign regs_120_reset = io_reset;
  assign regs_121_io_in = 64'h0;
  assign regs_121_io_init = 64'h0;
  assign regs_121_io_reset = reset;
  assign regs_121_io_enable = 1'h1;
  assign regs_121_clock = clock;
  assign regs_121_reset = io_reset;
  assign regs_122_io_in = 64'h0;
  assign regs_122_io_init = 64'h0;
  assign regs_122_io_reset = reset;
  assign regs_122_io_enable = 1'h1;
  assign regs_122_clock = clock;
  assign regs_122_reset = io_reset;
  assign regs_123_io_in = 64'h0;
  assign regs_123_io_init = 64'h0;
  assign regs_123_io_reset = reset;
  assign regs_123_io_enable = 1'h1;
  assign regs_123_clock = clock;
  assign regs_123_reset = io_reset;
  assign regs_124_io_in = 64'h0;
  assign regs_124_io_init = 64'h0;
  assign regs_124_io_reset = reset;
  assign regs_124_io_enable = 1'h1;
  assign regs_124_clock = clock;
  assign regs_124_reset = io_reset;
  assign regs_125_io_in = 64'h0;
  assign regs_125_io_init = 64'h0;
  assign regs_125_io_reset = reset;
  assign regs_125_io_enable = 1'h1;
  assign regs_125_clock = clock;
  assign regs_125_reset = io_reset;
  assign regs_126_io_in = 64'h0;
  assign regs_126_io_init = 64'h0;
  assign regs_126_io_reset = reset;
  assign regs_126_io_enable = 1'h1;
  assign regs_126_clock = clock;
  assign regs_126_reset = io_reset;
  assign regs_127_io_in = 64'h0;
  assign regs_127_io_init = 64'h0;
  assign regs_127_io_reset = reset;
  assign regs_127_io_enable = 1'h1;
  assign regs_127_clock = clock;
  assign regs_127_reset = io_reset;
  assign regs_128_io_in = 64'h0;
  assign regs_128_io_init = 64'h0;
  assign regs_128_io_reset = reset;
  assign regs_128_io_enable = 1'h1;
  assign regs_128_clock = clock;
  assign regs_128_reset = io_reset;
  assign regs_129_io_in = 64'h0;
  assign regs_129_io_init = 64'h0;
  assign regs_129_io_reset = reset;
  assign regs_129_io_enable = 1'h1;
  assign regs_129_clock = clock;
  assign regs_129_reset = io_reset;
  assign regs_130_io_in = 64'h0;
  assign regs_130_io_init = 64'h0;
  assign regs_130_io_reset = reset;
  assign regs_130_io_enable = 1'h1;
  assign regs_130_clock = clock;
  assign regs_130_reset = io_reset;
  assign regs_131_io_in = 64'h0;
  assign regs_131_io_init = 64'h0;
  assign regs_131_io_reset = reset;
  assign regs_131_io_enable = 1'h1;
  assign regs_131_clock = clock;
  assign regs_131_reset = io_reset;
  assign regs_132_io_in = 64'h0;
  assign regs_132_io_init = 64'h0;
  assign regs_132_io_reset = reset;
  assign regs_132_io_enable = 1'h1;
  assign regs_132_clock = clock;
  assign regs_132_reset = io_reset;
  assign regs_133_io_in = 64'h0;
  assign regs_133_io_init = 64'h0;
  assign regs_133_io_reset = reset;
  assign regs_133_io_enable = 1'h1;
  assign regs_133_clock = clock;
  assign regs_133_reset = io_reset;
  assign regs_134_io_in = 64'h0;
  assign regs_134_io_init = 64'h0;
  assign regs_134_io_reset = reset;
  assign regs_134_io_enable = 1'h1;
  assign regs_134_clock = clock;
  assign regs_134_reset = io_reset;
  assign regs_135_io_in = 64'h0;
  assign regs_135_io_init = 64'h0;
  assign regs_135_io_reset = reset;
  assign regs_135_io_enable = 1'h1;
  assign regs_135_clock = clock;
  assign regs_135_reset = io_reset;
  assign regs_136_io_in = 64'h0;
  assign regs_136_io_init = 64'h0;
  assign regs_136_io_reset = reset;
  assign regs_136_io_enable = 1'h1;
  assign regs_136_clock = clock;
  assign regs_136_reset = io_reset;
  assign regs_137_io_in = 64'h0;
  assign regs_137_io_init = 64'h0;
  assign regs_137_io_reset = reset;
  assign regs_137_io_enable = 1'h1;
  assign regs_137_clock = clock;
  assign regs_137_reset = io_reset;
  assign regs_138_io_in = 64'h0;
  assign regs_138_io_init = 64'h0;
  assign regs_138_io_reset = reset;
  assign regs_138_io_enable = 1'h1;
  assign regs_138_clock = clock;
  assign regs_138_reset = io_reset;
  assign regs_139_io_in = 64'h0;
  assign regs_139_io_init = 64'h0;
  assign regs_139_io_reset = reset;
  assign regs_139_io_enable = 1'h1;
  assign regs_139_clock = clock;
  assign regs_139_reset = io_reset;
  assign regs_140_io_in = 64'h0;
  assign regs_140_io_init = 64'h0;
  assign regs_140_io_reset = reset;
  assign regs_140_io_enable = 1'h1;
  assign regs_140_clock = clock;
  assign regs_140_reset = io_reset;
  assign regs_141_io_in = 64'h0;
  assign regs_141_io_init = 64'h0;
  assign regs_141_io_reset = reset;
  assign regs_141_io_enable = 1'h1;
  assign regs_141_clock = clock;
  assign regs_141_reset = io_reset;
  assign regs_142_io_in = 64'h0;
  assign regs_142_io_init = 64'h0;
  assign regs_142_io_reset = reset;
  assign regs_142_io_enable = 1'h1;
  assign regs_142_clock = clock;
  assign regs_142_reset = io_reset;
  assign regs_143_io_in = 64'h0;
  assign regs_143_io_init = 64'h0;
  assign regs_143_io_reset = reset;
  assign regs_143_io_enable = 1'h1;
  assign regs_143_clock = clock;
  assign regs_143_reset = io_reset;
  assign regs_144_io_in = 64'h0;
  assign regs_144_io_init = 64'h0;
  assign regs_144_io_reset = reset;
  assign regs_144_io_enable = 1'h1;
  assign regs_144_clock = clock;
  assign regs_144_reset = io_reset;
  assign regs_145_io_in = 64'h0;
  assign regs_145_io_init = 64'h0;
  assign regs_145_io_reset = reset;
  assign regs_145_io_enable = 1'h1;
  assign regs_145_clock = clock;
  assign regs_145_reset = io_reset;
  assign regs_146_io_in = 64'h0;
  assign regs_146_io_init = 64'h0;
  assign regs_146_io_reset = reset;
  assign regs_146_io_enable = 1'h1;
  assign regs_146_clock = clock;
  assign regs_146_reset = io_reset;
  assign regs_147_io_in = 64'h0;
  assign regs_147_io_init = 64'h0;
  assign regs_147_io_reset = reset;
  assign regs_147_io_enable = 1'h1;
  assign regs_147_clock = clock;
  assign regs_147_reset = io_reset;
  assign regs_148_io_in = 64'h0;
  assign regs_148_io_init = 64'h0;
  assign regs_148_io_reset = reset;
  assign regs_148_io_enable = 1'h1;
  assign regs_148_clock = clock;
  assign regs_148_reset = io_reset;
  assign regs_149_io_in = 64'h0;
  assign regs_149_io_init = 64'h0;
  assign regs_149_io_reset = reset;
  assign regs_149_io_enable = 1'h1;
  assign regs_149_clock = clock;
  assign regs_149_reset = io_reset;
  assign regs_150_io_in = 64'h0;
  assign regs_150_io_init = 64'h0;
  assign regs_150_io_reset = reset;
  assign regs_150_io_enable = 1'h1;
  assign regs_150_clock = clock;
  assign regs_150_reset = io_reset;
  assign regs_151_io_in = 64'h0;
  assign regs_151_io_init = 64'h0;
  assign regs_151_io_reset = reset;
  assign regs_151_io_enable = 1'h1;
  assign regs_151_clock = clock;
  assign regs_151_reset = io_reset;
  assign regs_152_io_in = 64'h0;
  assign regs_152_io_init = 64'h0;
  assign regs_152_io_reset = reset;
  assign regs_152_io_enable = 1'h1;
  assign regs_152_clock = clock;
  assign regs_152_reset = io_reset;
  assign regs_153_io_in = 64'h0;
  assign regs_153_io_init = 64'h0;
  assign regs_153_io_reset = reset;
  assign regs_153_io_enable = 1'h1;
  assign regs_153_clock = clock;
  assign regs_153_reset = io_reset;
  assign regs_154_io_in = 64'h0;
  assign regs_154_io_init = 64'h0;
  assign regs_154_io_reset = reset;
  assign regs_154_io_enable = 1'h1;
  assign regs_154_clock = clock;
  assign regs_154_reset = io_reset;
  assign regs_155_io_in = 64'h0;
  assign regs_155_io_init = 64'h0;
  assign regs_155_io_reset = reset;
  assign regs_155_io_enable = 1'h1;
  assign regs_155_clock = clock;
  assign regs_155_reset = io_reset;
  assign regs_156_io_in = 64'h0;
  assign regs_156_io_init = 64'h0;
  assign regs_156_io_reset = reset;
  assign regs_156_io_enable = 1'h1;
  assign regs_156_clock = clock;
  assign regs_156_reset = io_reset;
  assign regs_157_io_in = 64'h0;
  assign regs_157_io_init = 64'h0;
  assign regs_157_io_reset = reset;
  assign regs_157_io_enable = 1'h1;
  assign regs_157_clock = clock;
  assign regs_157_reset = io_reset;
  assign regs_158_io_in = 64'h0;
  assign regs_158_io_init = 64'h0;
  assign regs_158_io_reset = reset;
  assign regs_158_io_enable = 1'h1;
  assign regs_158_clock = clock;
  assign regs_158_reset = io_reset;
  assign regs_159_io_in = 64'h0;
  assign regs_159_io_init = 64'h0;
  assign regs_159_io_reset = reset;
  assign regs_159_io_enable = 1'h1;
  assign regs_159_clock = clock;
  assign regs_159_reset = io_reset;
  assign regs_160_io_in = 64'h0;
  assign regs_160_io_init = 64'h0;
  assign regs_160_io_reset = reset;
  assign regs_160_io_enable = 1'h1;
  assign regs_160_clock = clock;
  assign regs_160_reset = io_reset;
  assign regs_161_io_in = 64'h0;
  assign regs_161_io_init = 64'h0;
  assign regs_161_io_reset = reset;
  assign regs_161_io_enable = 1'h1;
  assign regs_161_clock = clock;
  assign regs_161_reset = io_reset;
  assign regs_162_io_in = 64'h0;
  assign regs_162_io_init = 64'h0;
  assign regs_162_io_reset = reset;
  assign regs_162_io_enable = 1'h1;
  assign regs_162_clock = clock;
  assign regs_162_reset = io_reset;
  assign regs_163_io_in = 64'h0;
  assign regs_163_io_init = 64'h0;
  assign regs_163_io_reset = reset;
  assign regs_163_io_enable = 1'h1;
  assign regs_163_clock = clock;
  assign regs_163_reset = io_reset;
  assign regs_164_io_in = 64'h0;
  assign regs_164_io_init = 64'h0;
  assign regs_164_io_reset = reset;
  assign regs_164_io_enable = 1'h1;
  assign regs_164_clock = clock;
  assign regs_164_reset = io_reset;
  assign regs_165_io_in = 64'h0;
  assign regs_165_io_init = 64'h0;
  assign regs_165_io_reset = reset;
  assign regs_165_io_enable = 1'h1;
  assign regs_165_clock = clock;
  assign regs_165_reset = io_reset;
  assign regs_166_io_in = 64'h0;
  assign regs_166_io_init = 64'h0;
  assign regs_166_io_reset = reset;
  assign regs_166_io_enable = 1'h1;
  assign regs_166_clock = clock;
  assign regs_166_reset = io_reset;
  assign regs_167_io_in = 64'h0;
  assign regs_167_io_init = 64'h0;
  assign regs_167_io_reset = reset;
  assign regs_167_io_enable = 1'h1;
  assign regs_167_clock = clock;
  assign regs_167_reset = io_reset;
  assign regs_168_io_in = 64'h0;
  assign regs_168_io_init = 64'h0;
  assign regs_168_io_reset = reset;
  assign regs_168_io_enable = 1'h1;
  assign regs_168_clock = clock;
  assign regs_168_reset = io_reset;
  assign regs_169_io_in = 64'h0;
  assign regs_169_io_init = 64'h0;
  assign regs_169_io_reset = reset;
  assign regs_169_io_enable = 1'h1;
  assign regs_169_clock = clock;
  assign regs_169_reset = io_reset;
  assign regs_170_io_in = 64'h0;
  assign regs_170_io_init = 64'h0;
  assign regs_170_io_reset = reset;
  assign regs_170_io_enable = 1'h1;
  assign regs_170_clock = clock;
  assign regs_170_reset = io_reset;
  assign regs_171_io_in = 64'h0;
  assign regs_171_io_init = 64'h0;
  assign regs_171_io_reset = reset;
  assign regs_171_io_enable = 1'h1;
  assign regs_171_clock = clock;
  assign regs_171_reset = io_reset;
  assign regs_172_io_in = 64'h0;
  assign regs_172_io_init = 64'h0;
  assign regs_172_io_reset = reset;
  assign regs_172_io_enable = 1'h1;
  assign regs_172_clock = clock;
  assign regs_172_reset = io_reset;
  assign regs_173_io_in = 64'h0;
  assign regs_173_io_init = 64'h0;
  assign regs_173_io_reset = reset;
  assign regs_173_io_enable = 1'h1;
  assign regs_173_clock = clock;
  assign regs_173_reset = io_reset;
  assign regs_174_io_in = 64'h0;
  assign regs_174_io_init = 64'h0;
  assign regs_174_io_reset = reset;
  assign regs_174_io_enable = 1'h1;
  assign regs_174_clock = clock;
  assign regs_174_reset = io_reset;
  assign regs_175_io_in = 64'h0;
  assign regs_175_io_init = 64'h0;
  assign regs_175_io_reset = reset;
  assign regs_175_io_enable = 1'h1;
  assign regs_175_clock = clock;
  assign regs_175_reset = io_reset;
  assign regs_176_io_in = 64'h0;
  assign regs_176_io_init = 64'h0;
  assign regs_176_io_reset = reset;
  assign regs_176_io_enable = 1'h1;
  assign regs_176_clock = clock;
  assign regs_176_reset = io_reset;
  assign regs_177_io_in = 64'h0;
  assign regs_177_io_init = 64'h0;
  assign regs_177_io_reset = reset;
  assign regs_177_io_enable = 1'h1;
  assign regs_177_clock = clock;
  assign regs_177_reset = io_reset;
  assign regs_178_io_in = 64'h0;
  assign regs_178_io_init = 64'h0;
  assign regs_178_io_reset = reset;
  assign regs_178_io_enable = 1'h1;
  assign regs_178_clock = clock;
  assign regs_178_reset = io_reset;
  assign regs_179_io_in = 64'h0;
  assign regs_179_io_init = 64'h0;
  assign regs_179_io_reset = reset;
  assign regs_179_io_enable = 1'h1;
  assign regs_179_clock = clock;
  assign regs_179_reset = io_reset;
  assign regs_180_io_in = 64'h0;
  assign regs_180_io_init = 64'h0;
  assign regs_180_io_reset = reset;
  assign regs_180_io_enable = 1'h1;
  assign regs_180_clock = clock;
  assign regs_180_reset = io_reset;
  assign regs_181_io_in = 64'h0;
  assign regs_181_io_init = 64'h0;
  assign regs_181_io_reset = reset;
  assign regs_181_io_enable = 1'h1;
  assign regs_181_clock = clock;
  assign regs_181_reset = io_reset;
  assign regs_182_io_in = 64'h0;
  assign regs_182_io_init = 64'h0;
  assign regs_182_io_reset = reset;
  assign regs_182_io_enable = 1'h1;
  assign regs_182_clock = clock;
  assign regs_182_reset = io_reset;
  assign regs_183_io_in = 64'h0;
  assign regs_183_io_init = 64'h0;
  assign regs_183_io_reset = reset;
  assign regs_183_io_enable = 1'h1;
  assign regs_183_clock = clock;
  assign regs_183_reset = io_reset;
  assign regs_184_io_in = 64'h0;
  assign regs_184_io_init = 64'h0;
  assign regs_184_io_reset = reset;
  assign regs_184_io_enable = 1'h1;
  assign regs_184_clock = clock;
  assign regs_184_reset = io_reset;
  assign regs_185_io_in = 64'h0;
  assign regs_185_io_init = 64'h0;
  assign regs_185_io_reset = reset;
  assign regs_185_io_enable = 1'h1;
  assign regs_185_clock = clock;
  assign regs_185_reset = io_reset;
  assign regs_186_io_in = 64'h0;
  assign regs_186_io_init = 64'h0;
  assign regs_186_io_reset = reset;
  assign regs_186_io_enable = 1'h1;
  assign regs_186_clock = clock;
  assign regs_186_reset = io_reset;
  assign regs_187_io_in = 64'h0;
  assign regs_187_io_init = 64'h0;
  assign regs_187_io_reset = reset;
  assign regs_187_io_enable = 1'h1;
  assign regs_187_clock = clock;
  assign regs_187_reset = io_reset;
  assign regs_188_io_in = 64'h0;
  assign regs_188_io_init = 64'h0;
  assign regs_188_io_reset = reset;
  assign regs_188_io_enable = 1'h1;
  assign regs_188_clock = clock;
  assign regs_188_reset = io_reset;
  assign regs_189_io_in = 64'h0;
  assign regs_189_io_init = 64'h0;
  assign regs_189_io_reset = reset;
  assign regs_189_io_enable = 1'h1;
  assign regs_189_clock = clock;
  assign regs_189_reset = io_reset;
  assign regs_190_io_in = 64'h0;
  assign regs_190_io_init = 64'h0;
  assign regs_190_io_reset = reset;
  assign regs_190_io_enable = 1'h1;
  assign regs_190_clock = clock;
  assign regs_190_reset = io_reset;
  assign regs_191_io_in = 64'h0;
  assign regs_191_io_init = 64'h0;
  assign regs_191_io_reset = reset;
  assign regs_191_io_enable = 1'h1;
  assign regs_191_clock = clock;
  assign regs_191_reset = io_reset;
  assign regs_192_io_in = 64'h0;
  assign regs_192_io_init = 64'h0;
  assign regs_192_io_reset = reset;
  assign regs_192_io_enable = 1'h1;
  assign regs_192_clock = clock;
  assign regs_192_reset = io_reset;
  assign regs_193_io_in = 64'h0;
  assign regs_193_io_init = 64'h0;
  assign regs_193_io_reset = reset;
  assign regs_193_io_enable = 1'h1;
  assign regs_193_clock = clock;
  assign regs_193_reset = io_reset;
  assign regs_194_io_in = 64'h0;
  assign regs_194_io_init = 64'h0;
  assign regs_194_io_reset = reset;
  assign regs_194_io_enable = 1'h1;
  assign regs_194_clock = clock;
  assign regs_194_reset = io_reset;
  assign regs_195_io_in = 64'h0;
  assign regs_195_io_init = 64'h0;
  assign regs_195_io_reset = reset;
  assign regs_195_io_enable = 1'h1;
  assign regs_195_clock = clock;
  assign regs_195_reset = io_reset;
  assign regs_196_io_in = 64'h0;
  assign regs_196_io_init = 64'h0;
  assign regs_196_io_reset = reset;
  assign regs_196_io_enable = 1'h1;
  assign regs_196_clock = clock;
  assign regs_196_reset = io_reset;
  assign regs_197_io_in = 64'h0;
  assign regs_197_io_init = 64'h0;
  assign regs_197_io_reset = reset;
  assign regs_197_io_enable = 1'h1;
  assign regs_197_clock = clock;
  assign regs_197_reset = io_reset;
  assign regs_198_io_in = 64'h0;
  assign regs_198_io_init = 64'h0;
  assign regs_198_io_reset = reset;
  assign regs_198_io_enable = 1'h1;
  assign regs_198_clock = clock;
  assign regs_198_reset = io_reset;
  assign regs_199_io_in = 64'h0;
  assign regs_199_io_init = 64'h0;
  assign regs_199_io_reset = reset;
  assign regs_199_io_enable = 1'h1;
  assign regs_199_clock = clock;
  assign regs_199_reset = io_reset;
  assign regs_200_io_in = 64'h0;
  assign regs_200_io_init = 64'h0;
  assign regs_200_io_reset = reset;
  assign regs_200_io_enable = 1'h1;
  assign regs_200_clock = clock;
  assign regs_200_reset = io_reset;
  assign regs_201_io_in = 64'h0;
  assign regs_201_io_init = 64'h0;
  assign regs_201_io_reset = reset;
  assign regs_201_io_enable = 1'h1;
  assign regs_201_clock = clock;
  assign regs_201_reset = io_reset;
  assign regs_202_io_in = 64'h0;
  assign regs_202_io_init = 64'h0;
  assign regs_202_io_reset = reset;
  assign regs_202_io_enable = 1'h1;
  assign regs_202_clock = clock;
  assign regs_202_reset = io_reset;
  assign regs_203_io_in = 64'h0;
  assign regs_203_io_init = 64'h0;
  assign regs_203_io_reset = reset;
  assign regs_203_io_enable = 1'h1;
  assign regs_203_clock = clock;
  assign regs_203_reset = io_reset;
  assign regs_204_io_in = 64'h0;
  assign regs_204_io_init = 64'h0;
  assign regs_204_io_reset = reset;
  assign regs_204_io_enable = 1'h1;
  assign regs_204_clock = clock;
  assign regs_204_reset = io_reset;
  assign regs_205_io_in = 64'h0;
  assign regs_205_io_init = 64'h0;
  assign regs_205_io_reset = reset;
  assign regs_205_io_enable = 1'h1;
  assign regs_205_clock = clock;
  assign regs_205_reset = io_reset;
  assign regs_206_io_in = 64'h0;
  assign regs_206_io_init = 64'h0;
  assign regs_206_io_reset = reset;
  assign regs_206_io_enable = 1'h1;
  assign regs_206_clock = clock;
  assign regs_206_reset = io_reset;
  assign regs_207_io_in = 64'h0;
  assign regs_207_io_init = 64'h0;
  assign regs_207_io_reset = reset;
  assign regs_207_io_enable = 1'h1;
  assign regs_207_clock = clock;
  assign regs_207_reset = io_reset;
  assign regs_208_io_in = 64'h0;
  assign regs_208_io_init = 64'h0;
  assign regs_208_io_reset = reset;
  assign regs_208_io_enable = 1'h1;
  assign regs_208_clock = clock;
  assign regs_208_reset = io_reset;
  assign regs_209_io_in = 64'h0;
  assign regs_209_io_init = 64'h0;
  assign regs_209_io_reset = reset;
  assign regs_209_io_enable = 1'h1;
  assign regs_209_clock = clock;
  assign regs_209_reset = io_reset;
  assign regs_210_io_in = 64'h0;
  assign regs_210_io_init = 64'h0;
  assign regs_210_io_reset = reset;
  assign regs_210_io_enable = 1'h1;
  assign regs_210_clock = clock;
  assign regs_210_reset = io_reset;
  assign regs_211_io_in = 64'h0;
  assign regs_211_io_init = 64'h0;
  assign regs_211_io_reset = reset;
  assign regs_211_io_enable = 1'h1;
  assign regs_211_clock = clock;
  assign regs_211_reset = io_reset;
  assign regs_212_io_in = 64'h0;
  assign regs_212_io_init = 64'h0;
  assign regs_212_io_reset = reset;
  assign regs_212_io_enable = 1'h1;
  assign regs_212_clock = clock;
  assign regs_212_reset = io_reset;
  assign regs_213_io_in = 64'h0;
  assign regs_213_io_init = 64'h0;
  assign regs_213_io_reset = reset;
  assign regs_213_io_enable = 1'h1;
  assign regs_213_clock = clock;
  assign regs_213_reset = io_reset;
  assign regs_214_io_in = 64'h0;
  assign regs_214_io_init = 64'h0;
  assign regs_214_io_reset = reset;
  assign regs_214_io_enable = 1'h1;
  assign regs_214_clock = clock;
  assign regs_214_reset = io_reset;
  assign regs_215_io_in = 64'h0;
  assign regs_215_io_init = 64'h0;
  assign regs_215_io_reset = reset;
  assign regs_215_io_enable = 1'h1;
  assign regs_215_clock = clock;
  assign regs_215_reset = io_reset;
  assign regs_216_io_in = 64'h0;
  assign regs_216_io_init = 64'h0;
  assign regs_216_io_reset = reset;
  assign regs_216_io_enable = 1'h1;
  assign regs_216_clock = clock;
  assign regs_216_reset = io_reset;
  assign regs_217_io_in = 64'h0;
  assign regs_217_io_init = 64'h0;
  assign regs_217_io_reset = reset;
  assign regs_217_io_enable = 1'h1;
  assign regs_217_clock = clock;
  assign regs_217_reset = io_reset;
  assign regs_218_io_in = 64'h0;
  assign regs_218_io_init = 64'h0;
  assign regs_218_io_reset = reset;
  assign regs_218_io_enable = 1'h1;
  assign regs_218_clock = clock;
  assign regs_218_reset = io_reset;
  assign regs_219_io_in = 64'h0;
  assign regs_219_io_init = 64'h0;
  assign regs_219_io_reset = reset;
  assign regs_219_io_enable = 1'h1;
  assign regs_219_clock = clock;
  assign regs_219_reset = io_reset;
  assign regs_220_io_in = 64'h0;
  assign regs_220_io_init = 64'h0;
  assign regs_220_io_reset = reset;
  assign regs_220_io_enable = 1'h1;
  assign regs_220_clock = clock;
  assign regs_220_reset = io_reset;
  assign regs_221_io_in = 64'h0;
  assign regs_221_io_init = 64'h0;
  assign regs_221_io_reset = reset;
  assign regs_221_io_enable = 1'h1;
  assign regs_221_clock = clock;
  assign regs_221_reset = io_reset;
  assign regs_222_io_in = 64'h0;
  assign regs_222_io_init = 64'h0;
  assign regs_222_io_reset = reset;
  assign regs_222_io_enable = 1'h1;
  assign regs_222_clock = clock;
  assign regs_222_reset = io_reset;
  assign regs_223_io_in = 64'h0;
  assign regs_223_io_init = 64'h0;
  assign regs_223_io_reset = reset;
  assign regs_223_io_enable = 1'h1;
  assign regs_223_clock = clock;
  assign regs_223_reset = io_reset;
  assign regs_224_io_in = 64'h0;
  assign regs_224_io_init = 64'h0;
  assign regs_224_io_reset = reset;
  assign regs_224_io_enable = 1'h1;
  assign regs_224_clock = clock;
  assign regs_224_reset = io_reset;
  assign regs_225_io_in = 64'h0;
  assign regs_225_io_init = 64'h0;
  assign regs_225_io_reset = reset;
  assign regs_225_io_enable = 1'h1;
  assign regs_225_clock = clock;
  assign regs_225_reset = io_reset;
  assign regs_226_io_in = 64'h0;
  assign regs_226_io_init = 64'h0;
  assign regs_226_io_reset = reset;
  assign regs_226_io_enable = 1'h1;
  assign regs_226_clock = clock;
  assign regs_226_reset = io_reset;
  assign regs_227_io_in = 64'h0;
  assign regs_227_io_init = 64'h0;
  assign regs_227_io_reset = reset;
  assign regs_227_io_enable = 1'h1;
  assign regs_227_clock = clock;
  assign regs_227_reset = io_reset;
  assign regs_228_io_in = 64'h0;
  assign regs_228_io_init = 64'h0;
  assign regs_228_io_reset = reset;
  assign regs_228_io_enable = 1'h1;
  assign regs_228_clock = clock;
  assign regs_228_reset = io_reset;
  assign regs_229_io_in = 64'h0;
  assign regs_229_io_init = 64'h0;
  assign regs_229_io_reset = reset;
  assign regs_229_io_enable = 1'h1;
  assign regs_229_clock = clock;
  assign regs_229_reset = io_reset;
  assign regs_230_io_in = 64'h0;
  assign regs_230_io_init = 64'h0;
  assign regs_230_io_reset = reset;
  assign regs_230_io_enable = 1'h1;
  assign regs_230_clock = clock;
  assign regs_230_reset = io_reset;
  assign regs_231_io_in = 64'h0;
  assign regs_231_io_init = 64'h0;
  assign regs_231_io_reset = reset;
  assign regs_231_io_enable = 1'h1;
  assign regs_231_clock = clock;
  assign regs_231_reset = io_reset;
  assign regs_232_io_in = 64'h0;
  assign regs_232_io_init = 64'h0;
  assign regs_232_io_reset = reset;
  assign regs_232_io_enable = 1'h1;
  assign regs_232_clock = clock;
  assign regs_232_reset = io_reset;
  assign regs_233_io_in = 64'h0;
  assign regs_233_io_init = 64'h0;
  assign regs_233_io_reset = reset;
  assign regs_233_io_enable = 1'h1;
  assign regs_233_clock = clock;
  assign regs_233_reset = io_reset;
  assign regs_234_io_in = 64'h0;
  assign regs_234_io_init = 64'h0;
  assign regs_234_io_reset = reset;
  assign regs_234_io_enable = 1'h1;
  assign regs_234_clock = clock;
  assign regs_234_reset = io_reset;
  assign regs_235_io_in = 64'h0;
  assign regs_235_io_init = 64'h0;
  assign regs_235_io_reset = reset;
  assign regs_235_io_enable = 1'h1;
  assign regs_235_clock = clock;
  assign regs_235_reset = io_reset;
  assign regs_236_io_in = 64'h0;
  assign regs_236_io_init = 64'h0;
  assign regs_236_io_reset = reset;
  assign regs_236_io_enable = 1'h1;
  assign regs_236_clock = clock;
  assign regs_236_reset = io_reset;
  assign regs_237_io_in = 64'h0;
  assign regs_237_io_init = 64'h0;
  assign regs_237_io_reset = reset;
  assign regs_237_io_enable = 1'h1;
  assign regs_237_clock = clock;
  assign regs_237_reset = io_reset;
  assign regs_238_io_in = 64'h0;
  assign regs_238_io_init = 64'h0;
  assign regs_238_io_reset = reset;
  assign regs_238_io_enable = 1'h1;
  assign regs_238_clock = clock;
  assign regs_238_reset = io_reset;
  assign regs_239_io_in = 64'h0;
  assign regs_239_io_init = 64'h0;
  assign regs_239_io_reset = reset;
  assign regs_239_io_enable = 1'h1;
  assign regs_239_clock = clock;
  assign regs_239_reset = io_reset;
  assign regs_240_io_in = 64'h0;
  assign regs_240_io_init = 64'h0;
  assign regs_240_io_reset = reset;
  assign regs_240_io_enable = 1'h1;
  assign regs_240_clock = clock;
  assign regs_240_reset = io_reset;
  assign regs_241_io_in = 64'h0;
  assign regs_241_io_init = 64'h0;
  assign regs_241_io_reset = reset;
  assign regs_241_io_enable = 1'h1;
  assign regs_241_clock = clock;
  assign regs_241_reset = io_reset;
  assign regs_242_io_in = 64'h0;
  assign regs_242_io_init = 64'h0;
  assign regs_242_io_reset = reset;
  assign regs_242_io_enable = 1'h1;
  assign regs_242_clock = clock;
  assign regs_242_reset = io_reset;
  assign regs_243_io_in = 64'h0;
  assign regs_243_io_init = 64'h0;
  assign regs_243_io_reset = reset;
  assign regs_243_io_enable = 1'h1;
  assign regs_243_clock = clock;
  assign regs_243_reset = io_reset;
  assign regs_244_io_in = 64'h0;
  assign regs_244_io_init = 64'h0;
  assign regs_244_io_reset = reset;
  assign regs_244_io_enable = 1'h1;
  assign regs_244_clock = clock;
  assign regs_244_reset = io_reset;
  assign regs_245_io_in = 64'h0;
  assign regs_245_io_init = 64'h0;
  assign regs_245_io_reset = reset;
  assign regs_245_io_enable = 1'h1;
  assign regs_245_clock = clock;
  assign regs_245_reset = io_reset;
  assign regs_246_io_in = 64'h0;
  assign regs_246_io_init = 64'h0;
  assign regs_246_io_reset = reset;
  assign regs_246_io_enable = 1'h1;
  assign regs_246_clock = clock;
  assign regs_246_reset = io_reset;
  assign regs_247_io_in = 64'h0;
  assign regs_247_io_init = 64'h0;
  assign regs_247_io_reset = reset;
  assign regs_247_io_enable = 1'h1;
  assign regs_247_clock = clock;
  assign regs_247_reset = io_reset;
  assign regs_248_io_in = 64'h0;
  assign regs_248_io_init = 64'h0;
  assign regs_248_io_reset = reset;
  assign regs_248_io_enable = 1'h1;
  assign regs_248_clock = clock;
  assign regs_248_reset = io_reset;
  assign regs_249_io_in = 64'h0;
  assign regs_249_io_init = 64'h0;
  assign regs_249_io_reset = reset;
  assign regs_249_io_enable = 1'h1;
  assign regs_249_clock = clock;
  assign regs_249_reset = io_reset;
  assign regs_250_io_in = 64'h0;
  assign regs_250_io_init = 64'h0;
  assign regs_250_io_reset = reset;
  assign regs_250_io_enable = 1'h1;
  assign regs_250_clock = clock;
  assign regs_250_reset = io_reset;
  assign regs_251_io_in = 64'h0;
  assign regs_251_io_init = 64'h0;
  assign regs_251_io_reset = reset;
  assign regs_251_io_enable = 1'h1;
  assign regs_251_clock = clock;
  assign regs_251_reset = io_reset;
  assign regs_252_io_in = 64'h0;
  assign regs_252_io_init = 64'h0;
  assign regs_252_io_reset = reset;
  assign regs_252_io_enable = 1'h1;
  assign regs_252_clock = clock;
  assign regs_252_reset = io_reset;
  assign regs_253_io_in = 64'h0;
  assign regs_253_io_init = 64'h0;
  assign regs_253_io_reset = reset;
  assign regs_253_io_enable = 1'h1;
  assign regs_253_clock = clock;
  assign regs_253_reset = io_reset;
  assign regs_254_io_in = 64'h0;
  assign regs_254_io_init = 64'h0;
  assign regs_254_io_reset = reset;
  assign regs_254_io_enable = 1'h1;
  assign regs_254_clock = clock;
  assign regs_254_reset = io_reset;
  assign regs_255_io_in = 64'h0;
  assign regs_255_io_init = 64'h0;
  assign regs_255_io_reset = reset;
  assign regs_255_io_enable = 1'h1;
  assign regs_255_clock = clock;
  assign regs_255_reset = io_reset;
  assign regs_256_io_in = 64'h0;
  assign regs_256_io_init = 64'h0;
  assign regs_256_io_reset = reset;
  assign regs_256_io_enable = 1'h1;
  assign regs_256_clock = clock;
  assign regs_256_reset = io_reset;
  assign regs_257_io_in = 64'h0;
  assign regs_257_io_init = 64'h0;
  assign regs_257_io_reset = reset;
  assign regs_257_io_enable = 1'h1;
  assign regs_257_clock = clock;
  assign regs_257_reset = io_reset;
  assign regs_258_io_in = 64'h0;
  assign regs_258_io_init = 64'h0;
  assign regs_258_io_reset = reset;
  assign regs_258_io_enable = 1'h1;
  assign regs_258_clock = clock;
  assign regs_258_reset = io_reset;
  assign regs_259_io_in = 64'h0;
  assign regs_259_io_init = 64'h0;
  assign regs_259_io_reset = reset;
  assign regs_259_io_enable = 1'h1;
  assign regs_259_clock = clock;
  assign regs_259_reset = io_reset;
  assign regs_260_io_in = 64'h0;
  assign regs_260_io_init = 64'h0;
  assign regs_260_io_reset = reset;
  assign regs_260_io_enable = 1'h1;
  assign regs_260_clock = clock;
  assign regs_260_reset = io_reset;
  assign regs_261_io_in = 64'h0;
  assign regs_261_io_init = 64'h0;
  assign regs_261_io_reset = reset;
  assign regs_261_io_enable = 1'h1;
  assign regs_261_clock = clock;
  assign regs_261_reset = io_reset;
  assign regs_262_io_in = 64'h0;
  assign regs_262_io_init = 64'h0;
  assign regs_262_io_reset = reset;
  assign regs_262_io_enable = 1'h1;
  assign regs_262_clock = clock;
  assign regs_262_reset = io_reset;
  assign regs_263_io_in = 64'h0;
  assign regs_263_io_init = 64'h0;
  assign regs_263_io_reset = reset;
  assign regs_263_io_enable = 1'h1;
  assign regs_263_clock = clock;
  assign regs_263_reset = io_reset;
  assign regs_264_io_in = 64'h0;
  assign regs_264_io_init = 64'h0;
  assign regs_264_io_reset = reset;
  assign regs_264_io_enable = 1'h1;
  assign regs_264_clock = clock;
  assign regs_264_reset = io_reset;
  assign regs_265_io_in = 64'h0;
  assign regs_265_io_init = 64'h0;
  assign regs_265_io_reset = reset;
  assign regs_265_io_enable = 1'h1;
  assign regs_265_clock = clock;
  assign regs_265_reset = io_reset;
  assign regs_266_io_in = 64'h0;
  assign regs_266_io_init = 64'h0;
  assign regs_266_io_reset = reset;
  assign regs_266_io_enable = 1'h1;
  assign regs_266_clock = clock;
  assign regs_266_reset = io_reset;
  assign regs_267_io_in = 64'h0;
  assign regs_267_io_init = 64'h0;
  assign regs_267_io_reset = reset;
  assign regs_267_io_enable = 1'h1;
  assign regs_267_clock = clock;
  assign regs_267_reset = io_reset;
  assign regs_268_io_in = 64'h0;
  assign regs_268_io_init = 64'h0;
  assign regs_268_io_reset = reset;
  assign regs_268_io_enable = 1'h1;
  assign regs_268_clock = clock;
  assign regs_268_reset = io_reset;
  assign regs_269_io_in = 64'h0;
  assign regs_269_io_init = 64'h0;
  assign regs_269_io_reset = reset;
  assign regs_269_io_enable = 1'h1;
  assign regs_269_clock = clock;
  assign regs_269_reset = io_reset;
  assign regs_270_io_in = 64'h0;
  assign regs_270_io_init = 64'h0;
  assign regs_270_io_reset = reset;
  assign regs_270_io_enable = 1'h1;
  assign regs_270_clock = clock;
  assign regs_270_reset = io_reset;
  assign regs_271_io_in = 64'h0;
  assign regs_271_io_init = 64'h0;
  assign regs_271_io_reset = reset;
  assign regs_271_io_enable = 1'h1;
  assign regs_271_clock = clock;
  assign regs_271_reset = io_reset;
  assign regs_272_io_in = 64'h0;
  assign regs_272_io_init = 64'h0;
  assign regs_272_io_reset = reset;
  assign regs_272_io_enable = 1'h1;
  assign regs_272_clock = clock;
  assign regs_272_reset = io_reset;
  assign regs_273_io_in = 64'h0;
  assign regs_273_io_init = 64'h0;
  assign regs_273_io_reset = reset;
  assign regs_273_io_enable = 1'h1;
  assign regs_273_clock = clock;
  assign regs_273_reset = io_reset;
  assign regs_274_io_in = 64'h0;
  assign regs_274_io_init = 64'h0;
  assign regs_274_io_reset = reset;
  assign regs_274_io_enable = 1'h1;
  assign regs_274_clock = clock;
  assign regs_274_reset = io_reset;
  assign regs_275_io_in = 64'h0;
  assign regs_275_io_init = 64'h0;
  assign regs_275_io_reset = reset;
  assign regs_275_io_enable = 1'h1;
  assign regs_275_clock = clock;
  assign regs_275_reset = io_reset;
  assign regs_276_io_in = 64'h0;
  assign regs_276_io_init = 64'h0;
  assign regs_276_io_reset = reset;
  assign regs_276_io_enable = 1'h1;
  assign regs_276_clock = clock;
  assign regs_276_reset = io_reset;
  assign regs_277_io_in = 64'h0;
  assign regs_277_io_init = 64'h0;
  assign regs_277_io_reset = reset;
  assign regs_277_io_enable = 1'h1;
  assign regs_277_clock = clock;
  assign regs_277_reset = io_reset;
  assign regs_278_io_in = 64'h0;
  assign regs_278_io_init = 64'h0;
  assign regs_278_io_reset = reset;
  assign regs_278_io_enable = 1'h1;
  assign regs_278_clock = clock;
  assign regs_278_reset = io_reset;
  assign regs_279_io_in = 64'h0;
  assign regs_279_io_init = 64'h0;
  assign regs_279_io_reset = reset;
  assign regs_279_io_enable = 1'h1;
  assign regs_279_clock = clock;
  assign regs_279_reset = io_reset;
  assign regs_280_io_in = 64'h0;
  assign regs_280_io_init = 64'h0;
  assign regs_280_io_reset = reset;
  assign regs_280_io_enable = 1'h1;
  assign regs_280_clock = clock;
  assign regs_280_reset = io_reset;
  assign regs_281_io_in = 64'h0;
  assign regs_281_io_init = 64'h0;
  assign regs_281_io_reset = reset;
  assign regs_281_io_enable = 1'h1;
  assign regs_281_clock = clock;
  assign regs_281_reset = io_reset;
  assign regs_282_io_in = 64'h0;
  assign regs_282_io_init = 64'h0;
  assign regs_282_io_reset = reset;
  assign regs_282_io_enable = 1'h1;
  assign regs_282_clock = clock;
  assign regs_282_reset = io_reset;
  assign regs_283_io_in = 64'h0;
  assign regs_283_io_init = 64'h0;
  assign regs_283_io_reset = reset;
  assign regs_283_io_enable = 1'h1;
  assign regs_283_clock = clock;
  assign regs_283_reset = io_reset;
  assign regs_284_io_in = 64'h0;
  assign regs_284_io_init = 64'h0;
  assign regs_284_io_reset = reset;
  assign regs_284_io_enable = 1'h1;
  assign regs_284_clock = clock;
  assign regs_284_reset = io_reset;
  assign regs_285_io_in = 64'h0;
  assign regs_285_io_init = 64'h0;
  assign regs_285_io_reset = reset;
  assign regs_285_io_enable = 1'h1;
  assign regs_285_clock = clock;
  assign regs_285_reset = io_reset;
  assign regs_286_io_in = 64'h0;
  assign regs_286_io_init = 64'h0;
  assign regs_286_io_reset = reset;
  assign regs_286_io_enable = 1'h1;
  assign regs_286_clock = clock;
  assign regs_286_reset = io_reset;
  assign regs_287_io_in = 64'h0;
  assign regs_287_io_init = 64'h0;
  assign regs_287_io_reset = reset;
  assign regs_287_io_enable = 1'h1;
  assign regs_287_clock = clock;
  assign regs_287_reset = io_reset;
  assign regs_288_io_in = 64'h0;
  assign regs_288_io_init = 64'h0;
  assign regs_288_io_reset = reset;
  assign regs_288_io_enable = 1'h1;
  assign regs_288_clock = clock;
  assign regs_288_reset = io_reset;
  assign regs_289_io_in = 64'h0;
  assign regs_289_io_init = 64'h0;
  assign regs_289_io_reset = reset;
  assign regs_289_io_enable = 1'h1;
  assign regs_289_clock = clock;
  assign regs_289_reset = io_reset;
  assign regs_290_io_in = 64'h0;
  assign regs_290_io_init = 64'h0;
  assign regs_290_io_reset = reset;
  assign regs_290_io_enable = 1'h1;
  assign regs_290_clock = clock;
  assign regs_290_reset = io_reset;
  assign regs_291_io_in = 64'h0;
  assign regs_291_io_init = 64'h0;
  assign regs_291_io_reset = reset;
  assign regs_291_io_enable = 1'h1;
  assign regs_291_clock = clock;
  assign regs_291_reset = io_reset;
  assign regs_292_io_in = 64'h0;
  assign regs_292_io_init = 64'h0;
  assign regs_292_io_reset = reset;
  assign regs_292_io_enable = 1'h1;
  assign regs_292_clock = clock;
  assign regs_292_reset = io_reset;
  assign regs_293_io_in = 64'h0;
  assign regs_293_io_init = 64'h0;
  assign regs_293_io_reset = reset;
  assign regs_293_io_enable = 1'h1;
  assign regs_293_clock = clock;
  assign regs_293_reset = io_reset;
  assign regs_294_io_in = 64'h0;
  assign regs_294_io_init = 64'h0;
  assign regs_294_io_reset = reset;
  assign regs_294_io_enable = 1'h1;
  assign regs_294_clock = clock;
  assign regs_294_reset = io_reset;
  assign regs_295_io_in = 64'h0;
  assign regs_295_io_init = 64'h0;
  assign regs_295_io_reset = reset;
  assign regs_295_io_enable = 1'h1;
  assign regs_295_clock = clock;
  assign regs_295_reset = io_reset;
  assign regs_296_io_in = 64'h0;
  assign regs_296_io_init = 64'h0;
  assign regs_296_io_reset = reset;
  assign regs_296_io_enable = 1'h1;
  assign regs_296_clock = clock;
  assign regs_296_reset = io_reset;
  assign regs_297_io_in = 64'h0;
  assign regs_297_io_init = 64'h0;
  assign regs_297_io_reset = reset;
  assign regs_297_io_enable = 1'h1;
  assign regs_297_clock = clock;
  assign regs_297_reset = io_reset;
  assign regs_298_io_in = 64'h0;
  assign regs_298_io_init = 64'h0;
  assign regs_298_io_reset = reset;
  assign regs_298_io_enable = 1'h1;
  assign regs_298_clock = clock;
  assign regs_298_reset = io_reset;
  assign regs_299_io_in = 64'h0;
  assign regs_299_io_init = 64'h0;
  assign regs_299_io_reset = reset;
  assign regs_299_io_enable = 1'h1;
  assign regs_299_clock = clock;
  assign regs_299_reset = io_reset;
  assign regs_300_io_in = 64'h0;
  assign regs_300_io_init = 64'h0;
  assign regs_300_io_reset = reset;
  assign regs_300_io_enable = 1'h1;
  assign regs_300_clock = clock;
  assign regs_300_reset = io_reset;
  assign regs_301_io_in = 64'h0;
  assign regs_301_io_init = 64'h0;
  assign regs_301_io_reset = reset;
  assign regs_301_io_enable = 1'h1;
  assign regs_301_clock = clock;
  assign regs_301_reset = io_reset;
  assign regs_302_io_in = 64'h0;
  assign regs_302_io_init = 64'h0;
  assign regs_302_io_reset = reset;
  assign regs_302_io_enable = 1'h1;
  assign regs_302_clock = clock;
  assign regs_302_reset = io_reset;
  assign regs_303_io_in = 64'h0;
  assign regs_303_io_init = 64'h0;
  assign regs_303_io_reset = reset;
  assign regs_303_io_enable = 1'h1;
  assign regs_303_clock = clock;
  assign regs_303_reset = io_reset;
  assign regs_304_io_in = 64'h0;
  assign regs_304_io_init = 64'h0;
  assign regs_304_io_reset = reset;
  assign regs_304_io_enable = 1'h1;
  assign regs_304_clock = clock;
  assign regs_304_reset = io_reset;
  assign regs_305_io_in = 64'h0;
  assign regs_305_io_init = 64'h0;
  assign regs_305_io_reset = reset;
  assign regs_305_io_enable = 1'h1;
  assign regs_305_clock = clock;
  assign regs_305_reset = io_reset;
  assign regs_306_io_in = 64'h0;
  assign regs_306_io_init = 64'h0;
  assign regs_306_io_reset = reset;
  assign regs_306_io_enable = 1'h1;
  assign regs_306_clock = clock;
  assign regs_306_reset = io_reset;
  assign regs_307_io_in = 64'h0;
  assign regs_307_io_init = 64'h0;
  assign regs_307_io_reset = reset;
  assign regs_307_io_enable = 1'h1;
  assign regs_307_clock = clock;
  assign regs_307_reset = io_reset;
  assign regs_308_io_in = 64'h0;
  assign regs_308_io_init = 64'h0;
  assign regs_308_io_reset = reset;
  assign regs_308_io_enable = 1'h1;
  assign regs_308_clock = clock;
  assign regs_308_reset = io_reset;
  assign regs_309_io_in = 64'h0;
  assign regs_309_io_init = 64'h0;
  assign regs_309_io_reset = reset;
  assign regs_309_io_enable = 1'h1;
  assign regs_309_clock = clock;
  assign regs_309_reset = io_reset;
  assign regs_310_io_in = 64'h0;
  assign regs_310_io_init = 64'h0;
  assign regs_310_io_reset = reset;
  assign regs_310_io_enable = 1'h1;
  assign regs_310_clock = clock;
  assign regs_310_reset = io_reset;
  assign regs_311_io_in = 64'h0;
  assign regs_311_io_init = 64'h0;
  assign regs_311_io_reset = reset;
  assign regs_311_io_enable = 1'h1;
  assign regs_311_clock = clock;
  assign regs_311_reset = io_reset;
  assign regs_312_io_in = 64'h0;
  assign regs_312_io_init = 64'h0;
  assign regs_312_io_reset = reset;
  assign regs_312_io_enable = 1'h1;
  assign regs_312_clock = clock;
  assign regs_312_reset = io_reset;
  assign regs_313_io_in = 64'h0;
  assign regs_313_io_init = 64'h0;
  assign regs_313_io_reset = reset;
  assign regs_313_io_enable = 1'h1;
  assign regs_313_clock = clock;
  assign regs_313_reset = io_reset;
  assign regs_314_io_in = 64'h0;
  assign regs_314_io_init = 64'h0;
  assign regs_314_io_reset = reset;
  assign regs_314_io_enable = 1'h1;
  assign regs_314_clock = clock;
  assign regs_314_reset = io_reset;
  assign regs_315_io_in = 64'h0;
  assign regs_315_io_init = 64'h0;
  assign regs_315_io_reset = reset;
  assign regs_315_io_enable = 1'h1;
  assign regs_315_clock = clock;
  assign regs_315_reset = io_reset;
  assign regs_316_io_in = 64'h0;
  assign regs_316_io_init = 64'h0;
  assign regs_316_io_reset = reset;
  assign regs_316_io_enable = 1'h1;
  assign regs_316_clock = clock;
  assign regs_316_reset = io_reset;
  assign regs_317_io_in = 64'h0;
  assign regs_317_io_init = 64'h0;
  assign regs_317_io_reset = reset;
  assign regs_317_io_enable = 1'h1;
  assign regs_317_clock = clock;
  assign regs_317_reset = io_reset;
  assign regs_318_io_in = 64'h0;
  assign regs_318_io_init = 64'h0;
  assign regs_318_io_reset = reset;
  assign regs_318_io_enable = 1'h1;
  assign regs_318_clock = clock;
  assign regs_318_reset = io_reset;
  assign regs_319_io_in = 64'h0;
  assign regs_319_io_init = 64'h0;
  assign regs_319_io_reset = reset;
  assign regs_319_io_enable = 1'h1;
  assign regs_319_clock = clock;
  assign regs_319_reset = io_reset;
  assign regs_320_io_in = 64'h0;
  assign regs_320_io_init = 64'h0;
  assign regs_320_io_reset = reset;
  assign regs_320_io_enable = 1'h1;
  assign regs_320_clock = clock;
  assign regs_320_reset = io_reset;
  assign regs_321_io_in = 64'h0;
  assign regs_321_io_init = 64'h0;
  assign regs_321_io_reset = reset;
  assign regs_321_io_enable = 1'h1;
  assign regs_321_clock = clock;
  assign regs_321_reset = io_reset;
  assign regs_322_io_in = 64'h0;
  assign regs_322_io_init = 64'h0;
  assign regs_322_io_reset = reset;
  assign regs_322_io_enable = 1'h1;
  assign regs_322_clock = clock;
  assign regs_322_reset = io_reset;
  assign regs_323_io_in = 64'h0;
  assign regs_323_io_init = 64'h0;
  assign regs_323_io_reset = reset;
  assign regs_323_io_enable = 1'h1;
  assign regs_323_clock = clock;
  assign regs_323_reset = io_reset;
  assign regs_324_io_in = 64'h0;
  assign regs_324_io_init = 64'h0;
  assign regs_324_io_reset = reset;
  assign regs_324_io_enable = 1'h1;
  assign regs_324_clock = clock;
  assign regs_324_reset = io_reset;
  assign regs_325_io_in = 64'h0;
  assign regs_325_io_init = 64'h0;
  assign regs_325_io_reset = reset;
  assign regs_325_io_enable = 1'h1;
  assign regs_325_clock = clock;
  assign regs_325_reset = io_reset;
  assign regs_326_io_in = 64'h0;
  assign regs_326_io_init = 64'h0;
  assign regs_326_io_reset = reset;
  assign regs_326_io_enable = 1'h1;
  assign regs_326_clock = clock;
  assign regs_326_reset = io_reset;
  assign regs_327_io_in = 64'h0;
  assign regs_327_io_init = 64'h0;
  assign regs_327_io_reset = reset;
  assign regs_327_io_enable = 1'h1;
  assign regs_327_clock = clock;
  assign regs_327_reset = io_reset;
  assign regs_328_io_in = 64'h0;
  assign regs_328_io_init = 64'h0;
  assign regs_328_io_reset = reset;
  assign regs_328_io_enable = 1'h1;
  assign regs_328_clock = clock;
  assign regs_328_reset = io_reset;
  assign regs_329_io_in = 64'h0;
  assign regs_329_io_init = 64'h0;
  assign regs_329_io_reset = reset;
  assign regs_329_io_enable = 1'h1;
  assign regs_329_clock = clock;
  assign regs_329_reset = io_reset;
  assign regs_330_io_in = 64'h0;
  assign regs_330_io_init = 64'h0;
  assign regs_330_io_reset = reset;
  assign regs_330_io_enable = 1'h1;
  assign regs_330_clock = clock;
  assign regs_330_reset = io_reset;
  assign regs_331_io_in = 64'h0;
  assign regs_331_io_init = 64'h0;
  assign regs_331_io_reset = reset;
  assign regs_331_io_enable = 1'h1;
  assign regs_331_clock = clock;
  assign regs_331_reset = io_reset;
  assign regs_332_io_in = 64'h0;
  assign regs_332_io_init = 64'h0;
  assign regs_332_io_reset = reset;
  assign regs_332_io_enable = 1'h1;
  assign regs_332_clock = clock;
  assign regs_332_reset = io_reset;
  assign regs_333_io_in = 64'h0;
  assign regs_333_io_init = 64'h0;
  assign regs_333_io_reset = reset;
  assign regs_333_io_enable = 1'h1;
  assign regs_333_clock = clock;
  assign regs_333_reset = io_reset;
  assign regs_334_io_in = 64'h0;
  assign regs_334_io_init = 64'h0;
  assign regs_334_io_reset = reset;
  assign regs_334_io_enable = 1'h1;
  assign regs_334_clock = clock;
  assign regs_334_reset = io_reset;
  assign regs_335_io_in = 64'h0;
  assign regs_335_io_init = 64'h0;
  assign regs_335_io_reset = reset;
  assign regs_335_io_enable = 1'h1;
  assign regs_335_clock = clock;
  assign regs_335_reset = io_reset;
  assign regs_336_io_in = 64'h0;
  assign regs_336_io_init = 64'h0;
  assign regs_336_io_reset = reset;
  assign regs_336_io_enable = 1'h1;
  assign regs_336_clock = clock;
  assign regs_336_reset = io_reset;
  assign regs_337_io_in = 64'h0;
  assign regs_337_io_init = 64'h0;
  assign regs_337_io_reset = reset;
  assign regs_337_io_enable = 1'h1;
  assign regs_337_clock = clock;
  assign regs_337_reset = io_reset;
  assign regs_338_io_in = 64'h0;
  assign regs_338_io_init = 64'h0;
  assign regs_338_io_reset = reset;
  assign regs_338_io_enable = 1'h1;
  assign regs_338_clock = clock;
  assign regs_338_reset = io_reset;
  assign regs_339_io_in = 64'h0;
  assign regs_339_io_init = 64'h0;
  assign regs_339_io_reset = reset;
  assign regs_339_io_enable = 1'h1;
  assign regs_339_clock = clock;
  assign regs_339_reset = io_reset;
  assign regs_340_io_in = 64'h0;
  assign regs_340_io_init = 64'h0;
  assign regs_340_io_reset = reset;
  assign regs_340_io_enable = 1'h1;
  assign regs_340_clock = clock;
  assign regs_340_reset = io_reset;
  assign regs_341_io_in = 64'h0;
  assign regs_341_io_init = 64'h0;
  assign regs_341_io_reset = reset;
  assign regs_341_io_enable = 1'h1;
  assign regs_341_clock = clock;
  assign regs_341_reset = io_reset;
  assign regs_342_io_in = 64'h0;
  assign regs_342_io_init = 64'h0;
  assign regs_342_io_reset = reset;
  assign regs_342_io_enable = 1'h1;
  assign regs_342_clock = clock;
  assign regs_342_reset = io_reset;
  assign regs_343_io_in = 64'h0;
  assign regs_343_io_init = 64'h0;
  assign regs_343_io_reset = reset;
  assign regs_343_io_enable = 1'h1;
  assign regs_343_clock = clock;
  assign regs_343_reset = io_reset;
  assign regs_344_io_in = 64'h0;
  assign regs_344_io_init = 64'h0;
  assign regs_344_io_reset = reset;
  assign regs_344_io_enable = 1'h1;
  assign regs_344_clock = clock;
  assign regs_344_reset = io_reset;
  assign regs_345_io_in = 64'h0;
  assign regs_345_io_init = 64'h0;
  assign regs_345_io_reset = reset;
  assign regs_345_io_enable = 1'h1;
  assign regs_345_clock = clock;
  assign regs_345_reset = io_reset;
  assign regs_346_io_in = 64'h0;
  assign regs_346_io_init = 64'h0;
  assign regs_346_io_reset = reset;
  assign regs_346_io_enable = 1'h1;
  assign regs_346_clock = clock;
  assign regs_346_reset = io_reset;
  assign regs_347_io_in = 64'h0;
  assign regs_347_io_init = 64'h0;
  assign regs_347_io_reset = reset;
  assign regs_347_io_enable = 1'h1;
  assign regs_347_clock = clock;
  assign regs_347_reset = io_reset;
  assign regs_348_io_in = 64'h0;
  assign regs_348_io_init = 64'h0;
  assign regs_348_io_reset = reset;
  assign regs_348_io_enable = 1'h1;
  assign regs_348_clock = clock;
  assign regs_348_reset = io_reset;
  assign regs_349_io_in = 64'h0;
  assign regs_349_io_init = 64'h0;
  assign regs_349_io_reset = reset;
  assign regs_349_io_enable = 1'h1;
  assign regs_349_clock = clock;
  assign regs_349_reset = io_reset;
  assign regs_350_io_in = 64'h0;
  assign regs_350_io_init = 64'h0;
  assign regs_350_io_reset = reset;
  assign regs_350_io_enable = 1'h1;
  assign regs_350_clock = clock;
  assign regs_350_reset = io_reset;
  assign regs_351_io_in = 64'h0;
  assign regs_351_io_init = 64'h0;
  assign regs_351_io_reset = reset;
  assign regs_351_io_enable = 1'h1;
  assign regs_351_clock = clock;
  assign regs_351_reset = io_reset;
  assign regs_352_io_in = 64'h0;
  assign regs_352_io_init = 64'h0;
  assign regs_352_io_reset = reset;
  assign regs_352_io_enable = 1'h1;
  assign regs_352_clock = clock;
  assign regs_352_reset = io_reset;
  assign regs_353_io_in = 64'h0;
  assign regs_353_io_init = 64'h0;
  assign regs_353_io_reset = reset;
  assign regs_353_io_enable = 1'h1;
  assign regs_353_clock = clock;
  assign regs_353_reset = io_reset;
  assign regs_354_io_in = 64'h0;
  assign regs_354_io_init = 64'h0;
  assign regs_354_io_reset = reset;
  assign regs_354_io_enable = 1'h1;
  assign regs_354_clock = clock;
  assign regs_354_reset = io_reset;
  assign regs_355_io_in = 64'h0;
  assign regs_355_io_init = 64'h0;
  assign regs_355_io_reset = reset;
  assign regs_355_io_enable = 1'h1;
  assign regs_355_clock = clock;
  assign regs_355_reset = io_reset;
  assign regs_356_io_in = 64'h0;
  assign regs_356_io_init = 64'h0;
  assign regs_356_io_reset = reset;
  assign regs_356_io_enable = 1'h1;
  assign regs_356_clock = clock;
  assign regs_356_reset = io_reset;
  assign regs_357_io_in = 64'h0;
  assign regs_357_io_init = 64'h0;
  assign regs_357_io_reset = reset;
  assign regs_357_io_enable = 1'h1;
  assign regs_357_clock = clock;
  assign regs_357_reset = io_reset;
  assign regs_358_io_in = 64'h0;
  assign regs_358_io_init = 64'h0;
  assign regs_358_io_reset = reset;
  assign regs_358_io_enable = 1'h1;
  assign regs_358_clock = clock;
  assign regs_358_reset = io_reset;
  assign regs_359_io_in = 64'h0;
  assign regs_359_io_init = 64'h0;
  assign regs_359_io_reset = reset;
  assign regs_359_io_enable = 1'h1;
  assign regs_359_clock = clock;
  assign regs_359_reset = io_reset;
  assign regs_360_io_in = 64'h0;
  assign regs_360_io_init = 64'h0;
  assign regs_360_io_reset = reset;
  assign regs_360_io_enable = 1'h1;
  assign regs_360_clock = clock;
  assign regs_360_reset = io_reset;
  assign regs_361_io_in = 64'h0;
  assign regs_361_io_init = 64'h0;
  assign regs_361_io_reset = reset;
  assign regs_361_io_enable = 1'h1;
  assign regs_361_clock = clock;
  assign regs_361_reset = io_reset;
  assign regs_362_io_in = 64'h0;
  assign regs_362_io_init = 64'h0;
  assign regs_362_io_reset = reset;
  assign regs_362_io_enable = 1'h1;
  assign regs_362_clock = clock;
  assign regs_362_reset = io_reset;
  assign regs_363_io_in = 64'h0;
  assign regs_363_io_init = 64'h0;
  assign regs_363_io_reset = reset;
  assign regs_363_io_enable = 1'h1;
  assign regs_363_clock = clock;
  assign regs_363_reset = io_reset;
  assign regs_364_io_in = 64'h0;
  assign regs_364_io_init = 64'h0;
  assign regs_364_io_reset = reset;
  assign regs_364_io_enable = 1'h1;
  assign regs_364_clock = clock;
  assign regs_364_reset = io_reset;
  assign regs_365_io_in = 64'h0;
  assign regs_365_io_init = 64'h0;
  assign regs_365_io_reset = reset;
  assign regs_365_io_enable = 1'h1;
  assign regs_365_clock = clock;
  assign regs_365_reset = io_reset;
  assign regs_366_io_in = 64'h0;
  assign regs_366_io_init = 64'h0;
  assign regs_366_io_reset = reset;
  assign regs_366_io_enable = 1'h1;
  assign regs_366_clock = clock;
  assign regs_366_reset = io_reset;
  assign regs_367_io_in = 64'h0;
  assign regs_367_io_init = 64'h0;
  assign regs_367_io_reset = reset;
  assign regs_367_io_enable = 1'h1;
  assign regs_367_clock = clock;
  assign regs_367_reset = io_reset;
  assign regs_368_io_in = 64'h0;
  assign regs_368_io_init = 64'h0;
  assign regs_368_io_reset = reset;
  assign regs_368_io_enable = 1'h1;
  assign regs_368_clock = clock;
  assign regs_368_reset = io_reset;
  assign regs_369_io_in = 64'h0;
  assign regs_369_io_init = 64'h0;
  assign regs_369_io_reset = reset;
  assign regs_369_io_enable = 1'h1;
  assign regs_369_clock = clock;
  assign regs_369_reset = io_reset;
  assign regs_370_io_in = 64'h0;
  assign regs_370_io_init = 64'h0;
  assign regs_370_io_reset = reset;
  assign regs_370_io_enable = 1'h1;
  assign regs_370_clock = clock;
  assign regs_370_reset = io_reset;
  assign regs_371_io_in = 64'h0;
  assign regs_371_io_init = 64'h0;
  assign regs_371_io_reset = reset;
  assign regs_371_io_enable = 1'h1;
  assign regs_371_clock = clock;
  assign regs_371_reset = io_reset;
  assign regs_372_io_in = 64'h0;
  assign regs_372_io_init = 64'h0;
  assign regs_372_io_reset = reset;
  assign regs_372_io_enable = 1'h1;
  assign regs_372_clock = clock;
  assign regs_372_reset = io_reset;
  assign regs_373_io_in = 64'h0;
  assign regs_373_io_init = 64'h0;
  assign regs_373_io_reset = reset;
  assign regs_373_io_enable = 1'h1;
  assign regs_373_clock = clock;
  assign regs_373_reset = io_reset;
  assign regs_374_io_in = 64'h0;
  assign regs_374_io_init = 64'h0;
  assign regs_374_io_reset = reset;
  assign regs_374_io_enable = 1'h1;
  assign regs_374_clock = clock;
  assign regs_374_reset = io_reset;
  assign regs_375_io_in = 64'h0;
  assign regs_375_io_init = 64'h0;
  assign regs_375_io_reset = reset;
  assign regs_375_io_enable = 1'h1;
  assign regs_375_clock = clock;
  assign regs_375_reset = io_reset;
  assign regs_376_io_in = 64'h0;
  assign regs_376_io_init = 64'h0;
  assign regs_376_io_reset = reset;
  assign regs_376_io_enable = 1'h1;
  assign regs_376_clock = clock;
  assign regs_376_reset = io_reset;
  assign regs_377_io_in = 64'h0;
  assign regs_377_io_init = 64'h0;
  assign regs_377_io_reset = reset;
  assign regs_377_io_enable = 1'h1;
  assign regs_377_clock = clock;
  assign regs_377_reset = io_reset;
  assign regs_378_io_in = 64'h0;
  assign regs_378_io_init = 64'h0;
  assign regs_378_io_reset = reset;
  assign regs_378_io_enable = 1'h1;
  assign regs_378_clock = clock;
  assign regs_378_reset = io_reset;
  assign regs_379_io_in = 64'h0;
  assign regs_379_io_init = 64'h0;
  assign regs_379_io_reset = reset;
  assign regs_379_io_enable = 1'h1;
  assign regs_379_clock = clock;
  assign regs_379_reset = io_reset;
  assign regs_380_io_in = 64'h0;
  assign regs_380_io_init = 64'h0;
  assign regs_380_io_reset = reset;
  assign regs_380_io_enable = 1'h1;
  assign regs_380_clock = clock;
  assign regs_380_reset = io_reset;
  assign regs_381_io_in = 64'h0;
  assign regs_381_io_init = 64'h0;
  assign regs_381_io_reset = reset;
  assign regs_381_io_enable = 1'h1;
  assign regs_381_clock = clock;
  assign regs_381_reset = io_reset;
  assign regs_382_io_in = 64'h0;
  assign regs_382_io_init = 64'h0;
  assign regs_382_io_reset = reset;
  assign regs_382_io_enable = 1'h1;
  assign regs_382_clock = clock;
  assign regs_382_reset = io_reset;
  assign regs_383_io_in = 64'h0;
  assign regs_383_io_init = 64'h0;
  assign regs_383_io_reset = reset;
  assign regs_383_io_enable = 1'h1;
  assign regs_383_clock = clock;
  assign regs_383_reset = io_reset;
  assign regs_384_io_in = 64'h0;
  assign regs_384_io_init = 64'h0;
  assign regs_384_io_reset = reset;
  assign regs_384_io_enable = 1'h1;
  assign regs_384_clock = clock;
  assign regs_384_reset = io_reset;
  assign regs_385_io_in = 64'h0;
  assign regs_385_io_init = 64'h0;
  assign regs_385_io_reset = reset;
  assign regs_385_io_enable = 1'h1;
  assign regs_385_clock = clock;
  assign regs_385_reset = io_reset;
  assign regs_386_io_in = 64'h0;
  assign regs_386_io_init = 64'h0;
  assign regs_386_io_reset = reset;
  assign regs_386_io_enable = 1'h1;
  assign regs_386_clock = clock;
  assign regs_386_reset = io_reset;
  assign regs_387_io_in = 64'h0;
  assign regs_387_io_init = 64'h0;
  assign regs_387_io_reset = reset;
  assign regs_387_io_enable = 1'h1;
  assign regs_387_clock = clock;
  assign regs_387_reset = io_reset;
  assign regs_388_io_in = 64'h0;
  assign regs_388_io_init = 64'h0;
  assign regs_388_io_reset = reset;
  assign regs_388_io_enable = 1'h1;
  assign regs_388_clock = clock;
  assign regs_388_reset = io_reset;
  assign regs_389_io_in = 64'h0;
  assign regs_389_io_init = 64'h0;
  assign regs_389_io_reset = reset;
  assign regs_389_io_enable = 1'h1;
  assign regs_389_clock = clock;
  assign regs_389_reset = io_reset;
  assign regs_390_io_in = 64'h0;
  assign regs_390_io_init = 64'h0;
  assign regs_390_io_reset = reset;
  assign regs_390_io_enable = 1'h1;
  assign regs_390_clock = clock;
  assign regs_390_reset = io_reset;
  assign regs_391_io_in = 64'h0;
  assign regs_391_io_init = 64'h0;
  assign regs_391_io_reset = reset;
  assign regs_391_io_enable = 1'h1;
  assign regs_391_clock = clock;
  assign regs_391_reset = io_reset;
  assign regs_392_io_in = 64'h0;
  assign regs_392_io_init = 64'h0;
  assign regs_392_io_reset = reset;
  assign regs_392_io_enable = 1'h1;
  assign regs_392_clock = clock;
  assign regs_392_reset = io_reset;
  assign regs_393_io_in = 64'h0;
  assign regs_393_io_init = 64'h0;
  assign regs_393_io_reset = reset;
  assign regs_393_io_enable = 1'h1;
  assign regs_393_clock = clock;
  assign regs_393_reset = io_reset;
  assign regs_394_io_in = 64'h0;
  assign regs_394_io_init = 64'h0;
  assign regs_394_io_reset = reset;
  assign regs_394_io_enable = 1'h1;
  assign regs_394_clock = clock;
  assign regs_394_reset = io_reset;
  assign regs_395_io_in = 64'h0;
  assign regs_395_io_init = 64'h0;
  assign regs_395_io_reset = reset;
  assign regs_395_io_enable = 1'h1;
  assign regs_395_clock = clock;
  assign regs_395_reset = io_reset;
  assign regs_396_io_in = 64'h0;
  assign regs_396_io_init = 64'h0;
  assign regs_396_io_reset = reset;
  assign regs_396_io_enable = 1'h1;
  assign regs_396_clock = clock;
  assign regs_396_reset = io_reset;
  assign regs_397_io_in = 64'h0;
  assign regs_397_io_init = 64'h0;
  assign regs_397_io_reset = reset;
  assign regs_397_io_enable = 1'h1;
  assign regs_397_clock = clock;
  assign regs_397_reset = io_reset;
  assign regs_398_io_in = 64'h0;
  assign regs_398_io_init = 64'h0;
  assign regs_398_io_reset = reset;
  assign regs_398_io_enable = 1'h1;
  assign regs_398_clock = clock;
  assign regs_398_reset = io_reset;
  assign regs_399_io_in = 64'h0;
  assign regs_399_io_init = 64'h0;
  assign regs_399_io_reset = reset;
  assign regs_399_io_enable = 1'h1;
  assign regs_399_clock = clock;
  assign regs_399_reset = io_reset;
  assign regs_400_io_in = 64'h0;
  assign regs_400_io_init = 64'h0;
  assign regs_400_io_reset = reset;
  assign regs_400_io_enable = 1'h1;
  assign regs_400_clock = clock;
  assign regs_400_reset = io_reset;
  assign regs_401_io_in = 64'h0;
  assign regs_401_io_init = 64'h0;
  assign regs_401_io_reset = reset;
  assign regs_401_io_enable = 1'h1;
  assign regs_401_clock = clock;
  assign regs_401_reset = io_reset;
  assign regs_402_io_in = 64'h0;
  assign regs_402_io_init = 64'h0;
  assign regs_402_io_reset = reset;
  assign regs_402_io_enable = 1'h1;
  assign regs_402_clock = clock;
  assign regs_402_reset = io_reset;
  assign regs_403_io_in = 64'h0;
  assign regs_403_io_init = 64'h0;
  assign regs_403_io_reset = reset;
  assign regs_403_io_enable = 1'h1;
  assign regs_403_clock = clock;
  assign regs_403_reset = io_reset;
  assign regs_404_io_in = 64'h0;
  assign regs_404_io_init = 64'h0;
  assign regs_404_io_reset = reset;
  assign regs_404_io_enable = 1'h1;
  assign regs_404_clock = clock;
  assign regs_404_reset = io_reset;
  assign regs_405_io_in = 64'h0;
  assign regs_405_io_init = 64'h0;
  assign regs_405_io_reset = reset;
  assign regs_405_io_enable = 1'h1;
  assign regs_405_clock = clock;
  assign regs_405_reset = io_reset;
  assign regs_406_io_in = 64'h0;
  assign regs_406_io_init = 64'h0;
  assign regs_406_io_reset = reset;
  assign regs_406_io_enable = 1'h1;
  assign regs_406_clock = clock;
  assign regs_406_reset = io_reset;
  assign regs_407_io_in = 64'h0;
  assign regs_407_io_init = 64'h0;
  assign regs_407_io_reset = reset;
  assign regs_407_io_enable = 1'h1;
  assign regs_407_clock = clock;
  assign regs_407_reset = io_reset;
  assign regs_408_io_in = 64'h0;
  assign regs_408_io_init = 64'h0;
  assign regs_408_io_reset = reset;
  assign regs_408_io_enable = 1'h1;
  assign regs_408_clock = clock;
  assign regs_408_reset = io_reset;
  assign regs_409_io_in = 64'h0;
  assign regs_409_io_init = 64'h0;
  assign regs_409_io_reset = reset;
  assign regs_409_io_enable = 1'h1;
  assign regs_409_clock = clock;
  assign regs_409_reset = io_reset;
  assign regs_410_io_in = 64'h0;
  assign regs_410_io_init = 64'h0;
  assign regs_410_io_reset = reset;
  assign regs_410_io_enable = 1'h1;
  assign regs_410_clock = clock;
  assign regs_410_reset = io_reset;
  assign regs_411_io_in = 64'h0;
  assign regs_411_io_init = 64'h0;
  assign regs_411_io_reset = reset;
  assign regs_411_io_enable = 1'h1;
  assign regs_411_clock = clock;
  assign regs_411_reset = io_reset;
  assign regs_412_io_in = 64'h0;
  assign regs_412_io_init = 64'h0;
  assign regs_412_io_reset = reset;
  assign regs_412_io_enable = 1'h1;
  assign regs_412_clock = clock;
  assign regs_412_reset = io_reset;
  assign regs_413_io_in = 64'h0;
  assign regs_413_io_init = 64'h0;
  assign regs_413_io_reset = reset;
  assign regs_413_io_enable = 1'h1;
  assign regs_413_clock = clock;
  assign regs_413_reset = io_reset;
  assign regs_414_io_in = 64'h0;
  assign regs_414_io_init = 64'h0;
  assign regs_414_io_reset = reset;
  assign regs_414_io_enable = 1'h1;
  assign regs_414_clock = clock;
  assign regs_414_reset = io_reset;
  assign regs_415_io_in = 64'h0;
  assign regs_415_io_init = 64'h0;
  assign regs_415_io_reset = reset;
  assign regs_415_io_enable = 1'h1;
  assign regs_415_clock = clock;
  assign regs_415_reset = io_reset;
  assign regs_416_io_in = 64'h0;
  assign regs_416_io_init = 64'h0;
  assign regs_416_io_reset = reset;
  assign regs_416_io_enable = 1'h1;
  assign regs_416_clock = clock;
  assign regs_416_reset = io_reset;
  assign regs_417_io_in = 64'h0;
  assign regs_417_io_init = 64'h0;
  assign regs_417_io_reset = reset;
  assign regs_417_io_enable = 1'h1;
  assign regs_417_clock = clock;
  assign regs_417_reset = io_reset;
  assign regs_418_io_in = 64'h0;
  assign regs_418_io_init = 64'h0;
  assign regs_418_io_reset = reset;
  assign regs_418_io_enable = 1'h1;
  assign regs_418_clock = clock;
  assign regs_418_reset = io_reset;
  assign regs_419_io_in = 64'h0;
  assign regs_419_io_init = 64'h0;
  assign regs_419_io_reset = reset;
  assign regs_419_io_enable = 1'h1;
  assign regs_419_clock = clock;
  assign regs_419_reset = io_reset;
  assign regs_420_io_in = 64'h0;
  assign regs_420_io_init = 64'h0;
  assign regs_420_io_reset = reset;
  assign regs_420_io_enable = 1'h1;
  assign regs_420_clock = clock;
  assign regs_420_reset = io_reset;
  assign regs_421_io_in = 64'h0;
  assign regs_421_io_init = 64'h0;
  assign regs_421_io_reset = reset;
  assign regs_421_io_enable = 1'h1;
  assign regs_421_clock = clock;
  assign regs_421_reset = io_reset;
  assign regs_422_io_in = 64'h0;
  assign regs_422_io_init = 64'h0;
  assign regs_422_io_reset = reset;
  assign regs_422_io_enable = 1'h1;
  assign regs_422_clock = clock;
  assign regs_422_reset = io_reset;
  assign regs_423_io_in = 64'h0;
  assign regs_423_io_init = 64'h0;
  assign regs_423_io_reset = reset;
  assign regs_423_io_enable = 1'h1;
  assign regs_423_clock = clock;
  assign regs_423_reset = io_reset;
  assign regs_424_io_in = 64'h0;
  assign regs_424_io_init = 64'h0;
  assign regs_424_io_reset = reset;
  assign regs_424_io_enable = 1'h1;
  assign regs_424_clock = clock;
  assign regs_424_reset = io_reset;
  assign regs_425_io_in = 64'h0;
  assign regs_425_io_init = 64'h0;
  assign regs_425_io_reset = reset;
  assign regs_425_io_enable = 1'h1;
  assign regs_425_clock = clock;
  assign regs_425_reset = io_reset;
  assign regs_426_io_in = 64'h0;
  assign regs_426_io_init = 64'h0;
  assign regs_426_io_reset = reset;
  assign regs_426_io_enable = 1'h1;
  assign regs_426_clock = clock;
  assign regs_426_reset = io_reset;
  assign regs_427_io_in = 64'h0;
  assign regs_427_io_init = 64'h0;
  assign regs_427_io_reset = reset;
  assign regs_427_io_enable = 1'h1;
  assign regs_427_clock = clock;
  assign regs_427_reset = io_reset;
  assign regs_428_io_in = 64'h0;
  assign regs_428_io_init = 64'h0;
  assign regs_428_io_reset = reset;
  assign regs_428_io_enable = 1'h1;
  assign regs_428_clock = clock;
  assign regs_428_reset = io_reset;
  assign regs_429_io_in = 64'h0;
  assign regs_429_io_init = 64'h0;
  assign regs_429_io_reset = reset;
  assign regs_429_io_enable = 1'h1;
  assign regs_429_clock = clock;
  assign regs_429_reset = io_reset;
  assign regs_430_io_in = 64'h0;
  assign regs_430_io_init = 64'h0;
  assign regs_430_io_reset = reset;
  assign regs_430_io_enable = 1'h1;
  assign regs_430_clock = clock;
  assign regs_430_reset = io_reset;
  assign regs_431_io_in = 64'h0;
  assign regs_431_io_init = 64'h0;
  assign regs_431_io_reset = reset;
  assign regs_431_io_enable = 1'h1;
  assign regs_431_clock = clock;
  assign regs_431_reset = io_reset;
  assign regs_432_io_in = 64'h0;
  assign regs_432_io_init = 64'h0;
  assign regs_432_io_reset = reset;
  assign regs_432_io_enable = 1'h1;
  assign regs_432_clock = clock;
  assign regs_432_reset = io_reset;
  assign regs_433_io_in = 64'h0;
  assign regs_433_io_init = 64'h0;
  assign regs_433_io_reset = reset;
  assign regs_433_io_enable = 1'h1;
  assign regs_433_clock = clock;
  assign regs_433_reset = io_reset;
  assign regs_434_io_in = 64'h0;
  assign regs_434_io_init = 64'h0;
  assign regs_434_io_reset = reset;
  assign regs_434_io_enable = 1'h1;
  assign regs_434_clock = clock;
  assign regs_434_reset = io_reset;
  assign regs_435_io_in = 64'h0;
  assign regs_435_io_init = 64'h0;
  assign regs_435_io_reset = reset;
  assign regs_435_io_enable = 1'h1;
  assign regs_435_clock = clock;
  assign regs_435_reset = io_reset;
  assign regs_436_io_in = 64'h0;
  assign regs_436_io_init = 64'h0;
  assign regs_436_io_reset = reset;
  assign regs_436_io_enable = 1'h1;
  assign regs_436_clock = clock;
  assign regs_436_reset = io_reset;
  assign regs_437_io_in = 64'h0;
  assign regs_437_io_init = 64'h0;
  assign regs_437_io_reset = reset;
  assign regs_437_io_enable = 1'h1;
  assign regs_437_clock = clock;
  assign regs_437_reset = io_reset;
  assign regs_438_io_in = 64'h0;
  assign regs_438_io_init = 64'h0;
  assign regs_438_io_reset = reset;
  assign regs_438_io_enable = 1'h1;
  assign regs_438_clock = clock;
  assign regs_438_reset = io_reset;
  assign regs_439_io_in = 64'h0;
  assign regs_439_io_init = 64'h0;
  assign regs_439_io_reset = reset;
  assign regs_439_io_enable = 1'h1;
  assign regs_439_clock = clock;
  assign regs_439_reset = io_reset;
  assign regs_440_io_in = 64'h0;
  assign regs_440_io_init = 64'h0;
  assign regs_440_io_reset = reset;
  assign regs_440_io_enable = 1'h1;
  assign regs_440_clock = clock;
  assign regs_440_reset = io_reset;
  assign regs_441_io_in = 64'h0;
  assign regs_441_io_init = 64'h0;
  assign regs_441_io_reset = reset;
  assign regs_441_io_enable = 1'h1;
  assign regs_441_clock = clock;
  assign regs_441_reset = io_reset;
  assign regs_442_io_in = 64'h0;
  assign regs_442_io_init = 64'h0;
  assign regs_442_io_reset = reset;
  assign regs_442_io_enable = 1'h1;
  assign regs_442_clock = clock;
  assign regs_442_reset = io_reset;
  assign regs_443_io_in = 64'h0;
  assign regs_443_io_init = 64'h0;
  assign regs_443_io_reset = reset;
  assign regs_443_io_enable = 1'h1;
  assign regs_443_clock = clock;
  assign regs_443_reset = io_reset;
  assign regs_444_io_in = 64'h0;
  assign regs_444_io_init = 64'h0;
  assign regs_444_io_reset = reset;
  assign regs_444_io_enable = 1'h1;
  assign regs_444_clock = clock;
  assign regs_444_reset = io_reset;
  assign regs_445_io_in = 64'h0;
  assign regs_445_io_init = 64'h0;
  assign regs_445_io_reset = reset;
  assign regs_445_io_enable = 1'h1;
  assign regs_445_clock = clock;
  assign regs_445_reset = io_reset;
  assign regs_446_io_in = 64'h0;
  assign regs_446_io_init = 64'h0;
  assign regs_446_io_reset = reset;
  assign regs_446_io_enable = 1'h1;
  assign regs_446_clock = clock;
  assign regs_446_reset = io_reset;
  assign regs_447_io_in = 64'h0;
  assign regs_447_io_init = 64'h0;
  assign regs_447_io_reset = reset;
  assign regs_447_io_enable = 1'h1;
  assign regs_447_clock = clock;
  assign regs_447_reset = io_reset;
  assign regs_448_io_in = 64'h0;
  assign regs_448_io_init = 64'h0;
  assign regs_448_io_reset = reset;
  assign regs_448_io_enable = 1'h1;
  assign regs_448_clock = clock;
  assign regs_448_reset = io_reset;
  assign regs_449_io_in = 64'h0;
  assign regs_449_io_init = 64'h0;
  assign regs_449_io_reset = reset;
  assign regs_449_io_enable = 1'h1;
  assign regs_449_clock = clock;
  assign regs_449_reset = io_reset;
  assign regs_450_io_in = 64'h0;
  assign regs_450_io_init = 64'h0;
  assign regs_450_io_reset = reset;
  assign regs_450_io_enable = 1'h1;
  assign regs_450_clock = clock;
  assign regs_450_reset = io_reset;
  assign regs_451_io_in = 64'h0;
  assign regs_451_io_init = 64'h0;
  assign regs_451_io_reset = reset;
  assign regs_451_io_enable = 1'h1;
  assign regs_451_clock = clock;
  assign regs_451_reset = io_reset;
  assign regs_452_io_in = 64'h0;
  assign regs_452_io_init = 64'h0;
  assign regs_452_io_reset = reset;
  assign regs_452_io_enable = 1'h1;
  assign regs_452_clock = clock;
  assign regs_452_reset = io_reset;
  assign regs_453_io_in = 64'h0;
  assign regs_453_io_init = 64'h0;
  assign regs_453_io_reset = reset;
  assign regs_453_io_enable = 1'h1;
  assign regs_453_clock = clock;
  assign regs_453_reset = io_reset;
  assign regs_454_io_in = 64'h0;
  assign regs_454_io_init = 64'h0;
  assign regs_454_io_reset = reset;
  assign regs_454_io_enable = 1'h1;
  assign regs_454_clock = clock;
  assign regs_454_reset = io_reset;
  assign regs_455_io_in = 64'h0;
  assign regs_455_io_init = 64'h0;
  assign regs_455_io_reset = reset;
  assign regs_455_io_enable = 1'h1;
  assign regs_455_clock = clock;
  assign regs_455_reset = io_reset;
  assign regs_456_io_in = 64'h0;
  assign regs_456_io_init = 64'h0;
  assign regs_456_io_reset = reset;
  assign regs_456_io_enable = 1'h1;
  assign regs_456_clock = clock;
  assign regs_456_reset = io_reset;
  assign regs_457_io_in = 64'h0;
  assign regs_457_io_init = 64'h0;
  assign regs_457_io_reset = reset;
  assign regs_457_io_enable = 1'h1;
  assign regs_457_clock = clock;
  assign regs_457_reset = io_reset;
  assign regs_458_io_in = 64'h0;
  assign regs_458_io_init = 64'h0;
  assign regs_458_io_reset = reset;
  assign regs_458_io_enable = 1'h1;
  assign regs_458_clock = clock;
  assign regs_458_reset = io_reset;
  assign regs_459_io_in = 64'h0;
  assign regs_459_io_init = 64'h0;
  assign regs_459_io_reset = reset;
  assign regs_459_io_enable = 1'h1;
  assign regs_459_clock = clock;
  assign regs_459_reset = io_reset;
  assign regs_460_io_in = 64'h0;
  assign regs_460_io_init = 64'h0;
  assign regs_460_io_reset = reset;
  assign regs_460_io_enable = 1'h1;
  assign regs_460_clock = clock;
  assign regs_460_reset = io_reset;
  assign regs_461_io_in = 64'h0;
  assign regs_461_io_init = 64'h0;
  assign regs_461_io_reset = reset;
  assign regs_461_io_enable = 1'h1;
  assign regs_461_clock = clock;
  assign regs_461_reset = io_reset;
  assign regs_462_io_in = 64'h0;
  assign regs_462_io_init = 64'h0;
  assign regs_462_io_reset = reset;
  assign regs_462_io_enable = 1'h1;
  assign regs_462_clock = clock;
  assign regs_462_reset = io_reset;
  assign regs_463_io_in = 64'h0;
  assign regs_463_io_init = 64'h0;
  assign regs_463_io_reset = reset;
  assign regs_463_io_enable = 1'h1;
  assign regs_463_clock = clock;
  assign regs_463_reset = io_reset;
  assign regs_464_io_in = 64'h0;
  assign regs_464_io_init = 64'h0;
  assign regs_464_io_reset = reset;
  assign regs_464_io_enable = 1'h1;
  assign regs_464_clock = clock;
  assign regs_464_reset = io_reset;
  assign regs_465_io_in = 64'h0;
  assign regs_465_io_init = 64'h0;
  assign regs_465_io_reset = reset;
  assign regs_465_io_enable = 1'h1;
  assign regs_465_clock = clock;
  assign regs_465_reset = io_reset;
  assign regs_466_io_in = 64'h0;
  assign regs_466_io_init = 64'h0;
  assign regs_466_io_reset = reset;
  assign regs_466_io_enable = 1'h1;
  assign regs_466_clock = clock;
  assign regs_466_reset = io_reset;
  assign regs_467_io_in = 64'h0;
  assign regs_467_io_init = 64'h0;
  assign regs_467_io_reset = reset;
  assign regs_467_io_enable = 1'h1;
  assign regs_467_clock = clock;
  assign regs_467_reset = io_reset;
  assign regs_468_io_in = 64'h0;
  assign regs_468_io_init = 64'h0;
  assign regs_468_io_reset = reset;
  assign regs_468_io_enable = 1'h1;
  assign regs_468_clock = clock;
  assign regs_468_reset = io_reset;
  assign regs_469_io_in = 64'h0;
  assign regs_469_io_init = 64'h0;
  assign regs_469_io_reset = reset;
  assign regs_469_io_enable = 1'h1;
  assign regs_469_clock = clock;
  assign regs_469_reset = io_reset;
  assign regs_470_io_in = 64'h0;
  assign regs_470_io_init = 64'h0;
  assign regs_470_io_reset = reset;
  assign regs_470_io_enable = 1'h1;
  assign regs_470_clock = clock;
  assign regs_470_reset = io_reset;
  assign regs_471_io_in = 64'h0;
  assign regs_471_io_init = 64'h0;
  assign regs_471_io_reset = reset;
  assign regs_471_io_enable = 1'h1;
  assign regs_471_clock = clock;
  assign regs_471_reset = io_reset;
  assign regs_472_io_in = 64'h0;
  assign regs_472_io_init = 64'h0;
  assign regs_472_io_reset = reset;
  assign regs_472_io_enable = 1'h1;
  assign regs_472_clock = clock;
  assign regs_472_reset = io_reset;
  assign regs_473_io_in = 64'h0;
  assign regs_473_io_init = 64'h0;
  assign regs_473_io_reset = reset;
  assign regs_473_io_enable = 1'h1;
  assign regs_473_clock = clock;
  assign regs_473_reset = io_reset;
  assign regs_474_io_in = 64'h0;
  assign regs_474_io_init = 64'h0;
  assign regs_474_io_reset = reset;
  assign regs_474_io_enable = 1'h1;
  assign regs_474_clock = clock;
  assign regs_474_reset = io_reset;
  assign regs_475_io_in = 64'h0;
  assign regs_475_io_init = 64'h0;
  assign regs_475_io_reset = reset;
  assign regs_475_io_enable = 1'h1;
  assign regs_475_clock = clock;
  assign regs_475_reset = io_reset;
  assign regs_476_io_in = 64'h0;
  assign regs_476_io_init = 64'h0;
  assign regs_476_io_reset = reset;
  assign regs_476_io_enable = 1'h1;
  assign regs_476_clock = clock;
  assign regs_476_reset = io_reset;
  assign regs_477_io_in = 64'h0;
  assign regs_477_io_init = 64'h0;
  assign regs_477_io_reset = reset;
  assign regs_477_io_enable = 1'h1;
  assign regs_477_clock = clock;
  assign regs_477_reset = io_reset;
  assign regs_478_io_in = 64'h0;
  assign regs_478_io_init = 64'h0;
  assign regs_478_io_reset = reset;
  assign regs_478_io_enable = 1'h1;
  assign regs_478_clock = clock;
  assign regs_478_reset = io_reset;
  assign regs_479_io_in = 64'h0;
  assign regs_479_io_init = 64'h0;
  assign regs_479_io_reset = reset;
  assign regs_479_io_enable = 1'h1;
  assign regs_479_clock = clock;
  assign regs_479_reset = io_reset;
  assign regs_480_io_in = 64'h0;
  assign regs_480_io_init = 64'h0;
  assign regs_480_io_reset = reset;
  assign regs_480_io_enable = 1'h1;
  assign regs_480_clock = clock;
  assign regs_480_reset = io_reset;
  assign regs_481_io_in = 64'h0;
  assign regs_481_io_init = 64'h0;
  assign regs_481_io_reset = reset;
  assign regs_481_io_enable = 1'h1;
  assign regs_481_clock = clock;
  assign regs_481_reset = io_reset;
  assign regs_482_io_in = 64'h0;
  assign regs_482_io_init = 64'h0;
  assign regs_482_io_reset = reset;
  assign regs_482_io_enable = 1'h1;
  assign regs_482_clock = clock;
  assign regs_482_reset = io_reset;
  assign regs_483_io_in = 64'h0;
  assign regs_483_io_init = 64'h0;
  assign regs_483_io_reset = reset;
  assign regs_483_io_enable = 1'h1;
  assign regs_483_clock = clock;
  assign regs_483_reset = io_reset;
  assign regs_484_io_in = 64'h0;
  assign regs_484_io_init = 64'h0;
  assign regs_484_io_reset = reset;
  assign regs_484_io_enable = 1'h1;
  assign regs_484_clock = clock;
  assign regs_484_reset = io_reset;
  assign regs_485_io_in = 64'h0;
  assign regs_485_io_init = 64'h0;
  assign regs_485_io_reset = reset;
  assign regs_485_io_enable = 1'h1;
  assign regs_485_clock = clock;
  assign regs_485_reset = io_reset;
  assign regs_486_io_in = 64'h0;
  assign regs_486_io_init = 64'h0;
  assign regs_486_io_reset = reset;
  assign regs_486_io_enable = 1'h1;
  assign regs_486_clock = clock;
  assign regs_486_reset = io_reset;
  assign regs_487_io_in = 64'h0;
  assign regs_487_io_init = 64'h0;
  assign regs_487_io_reset = reset;
  assign regs_487_io_enable = 1'h1;
  assign regs_487_clock = clock;
  assign regs_487_reset = io_reset;
  assign regs_488_io_in = 64'h0;
  assign regs_488_io_init = 64'h0;
  assign regs_488_io_reset = reset;
  assign regs_488_io_enable = 1'h1;
  assign regs_488_clock = clock;
  assign regs_488_reset = io_reset;
  assign regs_489_io_in = 64'h0;
  assign regs_489_io_init = 64'h0;
  assign regs_489_io_reset = reset;
  assign regs_489_io_enable = 1'h1;
  assign regs_489_clock = clock;
  assign regs_489_reset = io_reset;
  assign regs_490_io_in = 64'h0;
  assign regs_490_io_init = 64'h0;
  assign regs_490_io_reset = reset;
  assign regs_490_io_enable = 1'h1;
  assign regs_490_clock = clock;
  assign regs_490_reset = io_reset;
  assign regs_491_io_in = 64'h0;
  assign regs_491_io_init = 64'h0;
  assign regs_491_io_reset = reset;
  assign regs_491_io_enable = 1'h1;
  assign regs_491_clock = clock;
  assign regs_491_reset = io_reset;
  assign regs_492_io_in = 64'h0;
  assign regs_492_io_init = 64'h0;
  assign regs_492_io_reset = reset;
  assign regs_492_io_enable = 1'h1;
  assign regs_492_clock = clock;
  assign regs_492_reset = io_reset;
  assign regs_493_io_in = 64'h0;
  assign regs_493_io_init = 64'h0;
  assign regs_493_io_reset = reset;
  assign regs_493_io_enable = 1'h1;
  assign regs_493_clock = clock;
  assign regs_493_reset = io_reset;
  assign regs_494_io_in = 64'h0;
  assign regs_494_io_init = 64'h0;
  assign regs_494_io_reset = reset;
  assign regs_494_io_enable = 1'h1;
  assign regs_494_clock = clock;
  assign regs_494_reset = io_reset;
  assign regs_495_io_in = 64'h0;
  assign regs_495_io_init = 64'h0;
  assign regs_495_io_reset = reset;
  assign regs_495_io_enable = 1'h1;
  assign regs_495_clock = clock;
  assign regs_495_reset = io_reset;
  assign regs_496_io_in = 64'h0;
  assign regs_496_io_init = 64'h0;
  assign regs_496_io_reset = reset;
  assign regs_496_io_enable = 1'h1;
  assign regs_496_clock = clock;
  assign regs_496_reset = io_reset;
  assign regs_497_io_in = 64'h0;
  assign regs_497_io_init = 64'h0;
  assign regs_497_io_reset = reset;
  assign regs_497_io_enable = 1'h1;
  assign regs_497_clock = clock;
  assign regs_497_reset = io_reset;
  assign regs_498_io_in = 64'h0;
  assign regs_498_io_init = 64'h0;
  assign regs_498_io_reset = reset;
  assign regs_498_io_enable = 1'h1;
  assign regs_498_clock = clock;
  assign regs_498_reset = io_reset;
  assign regs_499_io_in = 64'h0;
  assign regs_499_io_init = 64'h0;
  assign regs_499_io_reset = reset;
  assign regs_499_io_enable = 1'h1;
  assign regs_499_clock = clock;
  assign regs_499_reset = io_reset;
  assign regs_500_io_in = 64'h0;
  assign regs_500_io_init = 64'h0;
  assign regs_500_io_reset = reset;
  assign regs_500_io_enable = 1'h1;
  assign regs_500_clock = clock;
  assign regs_500_reset = io_reset;
  assign regs_501_io_in = 64'h0;
  assign regs_501_io_init = 64'h0;
  assign regs_501_io_reset = reset;
  assign regs_501_io_enable = 1'h1;
  assign regs_501_clock = clock;
  assign regs_501_reset = io_reset;
  assign regs_502_io_in = 64'h0;
  assign regs_502_io_init = 64'h0;
  assign regs_502_io_reset = reset;
  assign regs_502_io_enable = 1'h1;
  assign regs_502_clock = clock;
  assign regs_502_reset = io_reset;
  assign regs_503_io_in = 64'h0;
  assign regs_503_io_init = 64'h0;
  assign regs_503_io_reset = reset;
  assign regs_503_io_enable = 1'h1;
  assign regs_503_clock = clock;
  assign regs_503_reset = io_reset;
  assign regs_504_io_in = 64'h0;
  assign regs_504_io_init = 64'h0;
  assign regs_504_io_reset = reset;
  assign regs_504_io_enable = 1'h1;
  assign regs_504_clock = clock;
  assign regs_504_reset = io_reset;
  assign regs_505_io_in = 64'h0;
  assign regs_505_io_init = 64'h0;
  assign regs_505_io_reset = reset;
  assign regs_505_io_enable = 1'h1;
  assign regs_505_clock = clock;
  assign regs_505_reset = io_reset;
  assign rport_io_ins_0 = regOuts_0;
  assign rport_io_ins_1 = regOuts_1;
  assign rport_io_ins_2 = regOuts_2;
  assign rport_io_ins_3 = regOuts_3;
  assign rport_io_ins_4 = regOuts_4;
  assign rport_io_ins_5 = regOuts_5;
  assign rport_io_ins_6 = regOuts_6;
  assign rport_io_ins_7 = regOuts_7;
  assign rport_io_ins_8 = regOuts_8;
  assign rport_io_ins_9 = regOuts_9;
  assign rport_io_ins_10 = regOuts_10;
  assign rport_io_ins_11 = regOuts_11;
  assign rport_io_ins_12 = regOuts_12;
  assign rport_io_ins_13 = regOuts_13;
  assign rport_io_ins_14 = regOuts_14;
  assign rport_io_ins_15 = regOuts_15;
  assign rport_io_ins_16 = regOuts_16;
  assign rport_io_ins_17 = regOuts_17;
  assign rport_io_ins_18 = regOuts_18;
  assign rport_io_ins_19 = regOuts_19;
  assign rport_io_ins_20 = regOuts_20;
  assign rport_io_ins_21 = regOuts_21;
  assign rport_io_ins_22 = regOuts_22;
  assign rport_io_ins_23 = regOuts_23;
  assign rport_io_ins_24 = regOuts_24;
  assign rport_io_ins_25 = regOuts_25;
  assign rport_io_ins_26 = regOuts_26;
  assign rport_io_ins_27 = regOuts_27;
  assign rport_io_ins_28 = regOuts_28;
  assign rport_io_ins_29 = regOuts_29;
  assign rport_io_ins_30 = regOuts_30;
  assign rport_io_ins_31 = regOuts_31;
  assign rport_io_ins_32 = regOuts_32;
  assign rport_io_ins_33 = regOuts_33;
  assign rport_io_ins_34 = regOuts_34;
  assign rport_io_ins_35 = regOuts_35;
  assign rport_io_ins_36 = regOuts_36;
  assign rport_io_ins_37 = regOuts_37;
  assign rport_io_ins_38 = regOuts_38;
  assign rport_io_ins_39 = regOuts_39;
  assign rport_io_ins_40 = regOuts_40;
  assign rport_io_ins_41 = regOuts_41;
  assign rport_io_ins_42 = regOuts_42;
  assign rport_io_ins_43 = regOuts_43;
  assign rport_io_ins_44 = regOuts_44;
  assign rport_io_ins_45 = regOuts_45;
  assign rport_io_ins_46 = regOuts_46;
  assign rport_io_ins_47 = regOuts_47;
  assign rport_io_ins_48 = regOuts_48;
  assign rport_io_ins_49 = regOuts_49;
  assign rport_io_ins_50 = regOuts_50;
  assign rport_io_ins_51 = regOuts_51;
  assign rport_io_ins_52 = regOuts_52;
  assign rport_io_ins_53 = regOuts_53;
  assign rport_io_ins_54 = regOuts_54;
  assign rport_io_ins_55 = regOuts_55;
  assign rport_io_ins_56 = regOuts_56;
  assign rport_io_ins_57 = regOuts_57;
  assign rport_io_ins_58 = regOuts_58;
  assign rport_io_ins_59 = regOuts_59;
  assign rport_io_ins_60 = regOuts_60;
  assign rport_io_ins_61 = regOuts_61;
  assign rport_io_ins_62 = regOuts_62;
  assign rport_io_ins_63 = regOuts_63;
  assign rport_io_ins_64 = regOuts_64;
  assign rport_io_ins_65 = regOuts_65;
  assign rport_io_ins_66 = regOuts_66;
  assign rport_io_ins_67 = regOuts_67;
  assign rport_io_ins_68 = regOuts_68;
  assign rport_io_ins_69 = regOuts_69;
  assign rport_io_ins_70 = regOuts_70;
  assign rport_io_ins_71 = regOuts_71;
  assign rport_io_ins_72 = regOuts_72;
  assign rport_io_ins_73 = regOuts_73;
  assign rport_io_ins_74 = regOuts_74;
  assign rport_io_ins_75 = regOuts_75;
  assign rport_io_ins_76 = regOuts_76;
  assign rport_io_ins_77 = regOuts_77;
  assign rport_io_ins_78 = regOuts_78;
  assign rport_io_ins_79 = regOuts_79;
  assign rport_io_ins_80 = regOuts_80;
  assign rport_io_ins_81 = regOuts_81;
  assign rport_io_ins_82 = regOuts_82;
  assign rport_io_ins_83 = regOuts_83;
  assign rport_io_ins_84 = regOuts_84;
  assign rport_io_ins_85 = regOuts_85;
  assign rport_io_ins_86 = regOuts_86;
  assign rport_io_ins_87 = regOuts_87;
  assign rport_io_ins_88 = regOuts_88;
  assign rport_io_ins_89 = regOuts_89;
  assign rport_io_ins_90 = regOuts_90;
  assign rport_io_ins_91 = regOuts_91;
  assign rport_io_ins_92 = regOuts_92;
  assign rport_io_ins_93 = regOuts_93;
  assign rport_io_ins_94 = regOuts_94;
  assign rport_io_ins_95 = regOuts_95;
  assign rport_io_ins_96 = regOuts_96;
  assign rport_io_ins_97 = regOuts_97;
  assign rport_io_ins_98 = regOuts_98;
  assign rport_io_ins_99 = regOuts_99;
  assign rport_io_ins_100 = regOuts_100;
  assign rport_io_ins_101 = regOuts_101;
  assign rport_io_ins_102 = regOuts_102;
  assign rport_io_ins_103 = regOuts_103;
  assign rport_io_ins_104 = regOuts_104;
  assign rport_io_ins_105 = regOuts_105;
  assign rport_io_ins_106 = regOuts_106;
  assign rport_io_ins_107 = regOuts_107;
  assign rport_io_ins_108 = regOuts_108;
  assign rport_io_ins_109 = regOuts_109;
  assign rport_io_ins_110 = regOuts_110;
  assign rport_io_ins_111 = regOuts_111;
  assign rport_io_ins_112 = regOuts_112;
  assign rport_io_ins_113 = regOuts_113;
  assign rport_io_ins_114 = regOuts_114;
  assign rport_io_ins_115 = regOuts_115;
  assign rport_io_ins_116 = regOuts_116;
  assign rport_io_ins_117 = regOuts_117;
  assign rport_io_ins_118 = regOuts_118;
  assign rport_io_ins_119 = regOuts_119;
  assign rport_io_ins_120 = regOuts_120;
  assign rport_io_ins_121 = regOuts_121;
  assign rport_io_ins_122 = regOuts_122;
  assign rport_io_ins_123 = regOuts_123;
  assign rport_io_ins_124 = regOuts_124;
  assign rport_io_ins_125 = regOuts_125;
  assign rport_io_ins_126 = regOuts_126;
  assign rport_io_ins_127 = regOuts_127;
  assign rport_io_ins_128 = regOuts_128;
  assign rport_io_ins_129 = regOuts_129;
  assign rport_io_ins_130 = regOuts_130;
  assign rport_io_ins_131 = regOuts_131;
  assign rport_io_ins_132 = regOuts_132;
  assign rport_io_ins_133 = regOuts_133;
  assign rport_io_ins_134 = regOuts_134;
  assign rport_io_ins_135 = regOuts_135;
  assign rport_io_ins_136 = regOuts_136;
  assign rport_io_ins_137 = regOuts_137;
  assign rport_io_ins_138 = regOuts_138;
  assign rport_io_ins_139 = regOuts_139;
  assign rport_io_ins_140 = regOuts_140;
  assign rport_io_ins_141 = regOuts_141;
  assign rport_io_ins_142 = regOuts_142;
  assign rport_io_ins_143 = regOuts_143;
  assign rport_io_ins_144 = regOuts_144;
  assign rport_io_ins_145 = regOuts_145;
  assign rport_io_ins_146 = regOuts_146;
  assign rport_io_ins_147 = regOuts_147;
  assign rport_io_ins_148 = regOuts_148;
  assign rport_io_ins_149 = regOuts_149;
  assign rport_io_ins_150 = regOuts_150;
  assign rport_io_ins_151 = regOuts_151;
  assign rport_io_ins_152 = regOuts_152;
  assign rport_io_ins_153 = regOuts_153;
  assign rport_io_ins_154 = regOuts_154;
  assign rport_io_ins_155 = regOuts_155;
  assign rport_io_ins_156 = regOuts_156;
  assign rport_io_ins_157 = regOuts_157;
  assign rport_io_ins_158 = regOuts_158;
  assign rport_io_ins_159 = regOuts_159;
  assign rport_io_ins_160 = regOuts_160;
  assign rport_io_ins_161 = regOuts_161;
  assign rport_io_ins_162 = regOuts_162;
  assign rport_io_ins_163 = regOuts_163;
  assign rport_io_ins_164 = regOuts_164;
  assign rport_io_ins_165 = regOuts_165;
  assign rport_io_ins_166 = regOuts_166;
  assign rport_io_ins_167 = regOuts_167;
  assign rport_io_ins_168 = regOuts_168;
  assign rport_io_ins_169 = regOuts_169;
  assign rport_io_ins_170 = regOuts_170;
  assign rport_io_ins_171 = regOuts_171;
  assign rport_io_ins_172 = regOuts_172;
  assign rport_io_ins_173 = regOuts_173;
  assign rport_io_ins_174 = regOuts_174;
  assign rport_io_ins_175 = regOuts_175;
  assign rport_io_ins_176 = regOuts_176;
  assign rport_io_ins_177 = regOuts_177;
  assign rport_io_ins_178 = regOuts_178;
  assign rport_io_ins_179 = regOuts_179;
  assign rport_io_ins_180 = regOuts_180;
  assign rport_io_ins_181 = regOuts_181;
  assign rport_io_ins_182 = regOuts_182;
  assign rport_io_ins_183 = regOuts_183;
  assign rport_io_ins_184 = regOuts_184;
  assign rport_io_ins_185 = regOuts_185;
  assign rport_io_ins_186 = regOuts_186;
  assign rport_io_ins_187 = regOuts_187;
  assign rport_io_ins_188 = regOuts_188;
  assign rport_io_ins_189 = regOuts_189;
  assign rport_io_ins_190 = regOuts_190;
  assign rport_io_ins_191 = regOuts_191;
  assign rport_io_ins_192 = regOuts_192;
  assign rport_io_ins_193 = regOuts_193;
  assign rport_io_ins_194 = regOuts_194;
  assign rport_io_ins_195 = regOuts_195;
  assign rport_io_ins_196 = regOuts_196;
  assign rport_io_ins_197 = regOuts_197;
  assign rport_io_ins_198 = regOuts_198;
  assign rport_io_ins_199 = regOuts_199;
  assign rport_io_ins_200 = regOuts_200;
  assign rport_io_ins_201 = regOuts_201;
  assign rport_io_ins_202 = regOuts_202;
  assign rport_io_ins_203 = regOuts_203;
  assign rport_io_ins_204 = regOuts_204;
  assign rport_io_ins_205 = regOuts_205;
  assign rport_io_ins_206 = regOuts_206;
  assign rport_io_ins_207 = regOuts_207;
  assign rport_io_ins_208 = regOuts_208;
  assign rport_io_ins_209 = regOuts_209;
  assign rport_io_ins_210 = regOuts_210;
  assign rport_io_ins_211 = regOuts_211;
  assign rport_io_ins_212 = regOuts_212;
  assign rport_io_ins_213 = regOuts_213;
  assign rport_io_ins_214 = regOuts_214;
  assign rport_io_ins_215 = regOuts_215;
  assign rport_io_ins_216 = regOuts_216;
  assign rport_io_ins_217 = regOuts_217;
  assign rport_io_ins_218 = regOuts_218;
  assign rport_io_ins_219 = regOuts_219;
  assign rport_io_ins_220 = regOuts_220;
  assign rport_io_ins_221 = regOuts_221;
  assign rport_io_ins_222 = regOuts_222;
  assign rport_io_ins_223 = regOuts_223;
  assign rport_io_ins_224 = regOuts_224;
  assign rport_io_ins_225 = regOuts_225;
  assign rport_io_ins_226 = regOuts_226;
  assign rport_io_ins_227 = regOuts_227;
  assign rport_io_ins_228 = regOuts_228;
  assign rport_io_ins_229 = regOuts_229;
  assign rport_io_ins_230 = regOuts_230;
  assign rport_io_ins_231 = regOuts_231;
  assign rport_io_ins_232 = regOuts_232;
  assign rport_io_ins_233 = regOuts_233;
  assign rport_io_ins_234 = regOuts_234;
  assign rport_io_ins_235 = regOuts_235;
  assign rport_io_ins_236 = regOuts_236;
  assign rport_io_ins_237 = regOuts_237;
  assign rport_io_ins_238 = regOuts_238;
  assign rport_io_ins_239 = regOuts_239;
  assign rport_io_ins_240 = regOuts_240;
  assign rport_io_ins_241 = regOuts_241;
  assign rport_io_ins_242 = regOuts_242;
  assign rport_io_ins_243 = regOuts_243;
  assign rport_io_ins_244 = regOuts_244;
  assign rport_io_ins_245 = regOuts_245;
  assign rport_io_ins_246 = regOuts_246;
  assign rport_io_ins_247 = regOuts_247;
  assign rport_io_ins_248 = regOuts_248;
  assign rport_io_ins_249 = regOuts_249;
  assign rport_io_ins_250 = regOuts_250;
  assign rport_io_ins_251 = regOuts_251;
  assign rport_io_ins_252 = regOuts_252;
  assign rport_io_ins_253 = regOuts_253;
  assign rport_io_ins_254 = regOuts_254;
  assign rport_io_ins_255 = regOuts_255;
  assign rport_io_ins_256 = regOuts_256;
  assign rport_io_ins_257 = regOuts_257;
  assign rport_io_ins_258 = regOuts_258;
  assign rport_io_ins_259 = regOuts_259;
  assign rport_io_ins_260 = regOuts_260;
  assign rport_io_ins_261 = regOuts_261;
  assign rport_io_ins_262 = regOuts_262;
  assign rport_io_ins_263 = regOuts_263;
  assign rport_io_ins_264 = regOuts_264;
  assign rport_io_ins_265 = regOuts_265;
  assign rport_io_ins_266 = regOuts_266;
  assign rport_io_ins_267 = regOuts_267;
  assign rport_io_ins_268 = regOuts_268;
  assign rport_io_ins_269 = regOuts_269;
  assign rport_io_ins_270 = regOuts_270;
  assign rport_io_ins_271 = regOuts_271;
  assign rport_io_ins_272 = regOuts_272;
  assign rport_io_ins_273 = regOuts_273;
  assign rport_io_ins_274 = regOuts_274;
  assign rport_io_ins_275 = regOuts_275;
  assign rport_io_ins_276 = regOuts_276;
  assign rport_io_ins_277 = regOuts_277;
  assign rport_io_ins_278 = regOuts_278;
  assign rport_io_ins_279 = regOuts_279;
  assign rport_io_ins_280 = regOuts_280;
  assign rport_io_ins_281 = regOuts_281;
  assign rport_io_ins_282 = regOuts_282;
  assign rport_io_ins_283 = regOuts_283;
  assign rport_io_ins_284 = regOuts_284;
  assign rport_io_ins_285 = regOuts_285;
  assign rport_io_ins_286 = regOuts_286;
  assign rport_io_ins_287 = regOuts_287;
  assign rport_io_ins_288 = regOuts_288;
  assign rport_io_ins_289 = regOuts_289;
  assign rport_io_ins_290 = regOuts_290;
  assign rport_io_ins_291 = regOuts_291;
  assign rport_io_ins_292 = regOuts_292;
  assign rport_io_ins_293 = regOuts_293;
  assign rport_io_ins_294 = regOuts_294;
  assign rport_io_ins_295 = regOuts_295;
  assign rport_io_ins_296 = regOuts_296;
  assign rport_io_ins_297 = regOuts_297;
  assign rport_io_ins_298 = regOuts_298;
  assign rport_io_ins_299 = regOuts_299;
  assign rport_io_ins_300 = regOuts_300;
  assign rport_io_ins_301 = regOuts_301;
  assign rport_io_ins_302 = regOuts_302;
  assign rport_io_ins_303 = regOuts_303;
  assign rport_io_ins_304 = regOuts_304;
  assign rport_io_ins_305 = regOuts_305;
  assign rport_io_ins_306 = regOuts_306;
  assign rport_io_ins_307 = regOuts_307;
  assign rport_io_ins_308 = regOuts_308;
  assign rport_io_ins_309 = regOuts_309;
  assign rport_io_ins_310 = regOuts_310;
  assign rport_io_ins_311 = regOuts_311;
  assign rport_io_ins_312 = regOuts_312;
  assign rport_io_ins_313 = regOuts_313;
  assign rport_io_ins_314 = regOuts_314;
  assign rport_io_ins_315 = regOuts_315;
  assign rport_io_ins_316 = regOuts_316;
  assign rport_io_ins_317 = regOuts_317;
  assign rport_io_ins_318 = regOuts_318;
  assign rport_io_ins_319 = regOuts_319;
  assign rport_io_ins_320 = regOuts_320;
  assign rport_io_ins_321 = regOuts_321;
  assign rport_io_ins_322 = regOuts_322;
  assign rport_io_ins_323 = regOuts_323;
  assign rport_io_ins_324 = regOuts_324;
  assign rport_io_ins_325 = regOuts_325;
  assign rport_io_ins_326 = regOuts_326;
  assign rport_io_ins_327 = regOuts_327;
  assign rport_io_ins_328 = regOuts_328;
  assign rport_io_ins_329 = regOuts_329;
  assign rport_io_ins_330 = regOuts_330;
  assign rport_io_ins_331 = regOuts_331;
  assign rport_io_ins_332 = regOuts_332;
  assign rport_io_ins_333 = regOuts_333;
  assign rport_io_ins_334 = regOuts_334;
  assign rport_io_ins_335 = regOuts_335;
  assign rport_io_ins_336 = regOuts_336;
  assign rport_io_ins_337 = regOuts_337;
  assign rport_io_ins_338 = regOuts_338;
  assign rport_io_ins_339 = regOuts_339;
  assign rport_io_ins_340 = regOuts_340;
  assign rport_io_ins_341 = regOuts_341;
  assign rport_io_ins_342 = regOuts_342;
  assign rport_io_ins_343 = regOuts_343;
  assign rport_io_ins_344 = regOuts_344;
  assign rport_io_ins_345 = regOuts_345;
  assign rport_io_ins_346 = regOuts_346;
  assign rport_io_ins_347 = regOuts_347;
  assign rport_io_ins_348 = regOuts_348;
  assign rport_io_ins_349 = regOuts_349;
  assign rport_io_ins_350 = regOuts_350;
  assign rport_io_ins_351 = regOuts_351;
  assign rport_io_ins_352 = regOuts_352;
  assign rport_io_ins_353 = regOuts_353;
  assign rport_io_ins_354 = regOuts_354;
  assign rport_io_ins_355 = regOuts_355;
  assign rport_io_ins_356 = regOuts_356;
  assign rport_io_ins_357 = regOuts_357;
  assign rport_io_ins_358 = regOuts_358;
  assign rport_io_ins_359 = regOuts_359;
  assign rport_io_ins_360 = regOuts_360;
  assign rport_io_ins_361 = regOuts_361;
  assign rport_io_ins_362 = regOuts_362;
  assign rport_io_ins_363 = regOuts_363;
  assign rport_io_ins_364 = regOuts_364;
  assign rport_io_ins_365 = regOuts_365;
  assign rport_io_ins_366 = regOuts_366;
  assign rport_io_ins_367 = regOuts_367;
  assign rport_io_ins_368 = regOuts_368;
  assign rport_io_ins_369 = regOuts_369;
  assign rport_io_ins_370 = regOuts_370;
  assign rport_io_ins_371 = regOuts_371;
  assign rport_io_ins_372 = regOuts_372;
  assign rport_io_ins_373 = regOuts_373;
  assign rport_io_ins_374 = regOuts_374;
  assign rport_io_ins_375 = regOuts_375;
  assign rport_io_ins_376 = regOuts_376;
  assign rport_io_ins_377 = regOuts_377;
  assign rport_io_ins_378 = regOuts_378;
  assign rport_io_ins_379 = regOuts_379;
  assign rport_io_ins_380 = regOuts_380;
  assign rport_io_ins_381 = regOuts_381;
  assign rport_io_ins_382 = regOuts_382;
  assign rport_io_ins_383 = regOuts_383;
  assign rport_io_ins_384 = regOuts_384;
  assign rport_io_ins_385 = regOuts_385;
  assign rport_io_ins_386 = regOuts_386;
  assign rport_io_ins_387 = regOuts_387;
  assign rport_io_ins_388 = regOuts_388;
  assign rport_io_ins_389 = regOuts_389;
  assign rport_io_ins_390 = regOuts_390;
  assign rport_io_ins_391 = regOuts_391;
  assign rport_io_ins_392 = regOuts_392;
  assign rport_io_ins_393 = regOuts_393;
  assign rport_io_ins_394 = regOuts_394;
  assign rport_io_ins_395 = regOuts_395;
  assign rport_io_ins_396 = regOuts_396;
  assign rport_io_ins_397 = regOuts_397;
  assign rport_io_ins_398 = regOuts_398;
  assign rport_io_ins_399 = regOuts_399;
  assign rport_io_ins_400 = regOuts_400;
  assign rport_io_ins_401 = regOuts_401;
  assign rport_io_ins_402 = regOuts_402;
  assign rport_io_ins_403 = regOuts_403;
  assign rport_io_ins_404 = regOuts_404;
  assign rport_io_ins_405 = regOuts_405;
  assign rport_io_ins_406 = regOuts_406;
  assign rport_io_ins_407 = regOuts_407;
  assign rport_io_ins_408 = regOuts_408;
  assign rport_io_ins_409 = regOuts_409;
  assign rport_io_ins_410 = regOuts_410;
  assign rport_io_ins_411 = regOuts_411;
  assign rport_io_ins_412 = regOuts_412;
  assign rport_io_ins_413 = regOuts_413;
  assign rport_io_ins_414 = regOuts_414;
  assign rport_io_ins_415 = regOuts_415;
  assign rport_io_ins_416 = regOuts_416;
  assign rport_io_ins_417 = regOuts_417;
  assign rport_io_ins_418 = regOuts_418;
  assign rport_io_ins_419 = regOuts_419;
  assign rport_io_ins_420 = regOuts_420;
  assign rport_io_ins_421 = regOuts_421;
  assign rport_io_ins_422 = regOuts_422;
  assign rport_io_ins_423 = regOuts_423;
  assign rport_io_ins_424 = regOuts_424;
  assign rport_io_ins_425 = regOuts_425;
  assign rport_io_ins_426 = regOuts_426;
  assign rport_io_ins_427 = regOuts_427;
  assign rport_io_ins_428 = regOuts_428;
  assign rport_io_ins_429 = regOuts_429;
  assign rport_io_ins_430 = regOuts_430;
  assign rport_io_ins_431 = regOuts_431;
  assign rport_io_ins_432 = regOuts_432;
  assign rport_io_ins_433 = regOuts_433;
  assign rport_io_ins_434 = regOuts_434;
  assign rport_io_ins_435 = regOuts_435;
  assign rport_io_ins_436 = regOuts_436;
  assign rport_io_ins_437 = regOuts_437;
  assign rport_io_ins_438 = regOuts_438;
  assign rport_io_ins_439 = regOuts_439;
  assign rport_io_ins_440 = regOuts_440;
  assign rport_io_ins_441 = regOuts_441;
  assign rport_io_ins_442 = regOuts_442;
  assign rport_io_ins_443 = regOuts_443;
  assign rport_io_ins_444 = regOuts_444;
  assign rport_io_ins_445 = regOuts_445;
  assign rport_io_ins_446 = regOuts_446;
  assign rport_io_ins_447 = regOuts_447;
  assign rport_io_ins_448 = regOuts_448;
  assign rport_io_ins_449 = regOuts_449;
  assign rport_io_ins_450 = regOuts_450;
  assign rport_io_ins_451 = regOuts_451;
  assign rport_io_ins_452 = regOuts_452;
  assign rport_io_ins_453 = regOuts_453;
  assign rport_io_ins_454 = regOuts_454;
  assign rport_io_ins_455 = regOuts_455;
  assign rport_io_ins_456 = regOuts_456;
  assign rport_io_ins_457 = regOuts_457;
  assign rport_io_ins_458 = regOuts_458;
  assign rport_io_ins_459 = regOuts_459;
  assign rport_io_ins_460 = regOuts_460;
  assign rport_io_ins_461 = regOuts_461;
  assign rport_io_ins_462 = regOuts_462;
  assign rport_io_ins_463 = regOuts_463;
  assign rport_io_ins_464 = regOuts_464;
  assign rport_io_ins_465 = regOuts_465;
  assign rport_io_ins_466 = regOuts_466;
  assign rport_io_ins_467 = regOuts_467;
  assign rport_io_ins_468 = regOuts_468;
  assign rport_io_ins_469 = regOuts_469;
  assign rport_io_ins_470 = regOuts_470;
  assign rport_io_ins_471 = regOuts_471;
  assign rport_io_ins_472 = regOuts_472;
  assign rport_io_ins_473 = regOuts_473;
  assign rport_io_ins_474 = regOuts_474;
  assign rport_io_ins_475 = regOuts_475;
  assign rport_io_ins_476 = regOuts_476;
  assign rport_io_ins_477 = regOuts_477;
  assign rport_io_ins_478 = regOuts_478;
  assign rport_io_ins_479 = regOuts_479;
  assign rport_io_ins_480 = regOuts_480;
  assign rport_io_ins_481 = regOuts_481;
  assign rport_io_ins_482 = regOuts_482;
  assign rport_io_ins_483 = regOuts_483;
  assign rport_io_ins_484 = regOuts_484;
  assign rport_io_ins_485 = regOuts_485;
  assign rport_io_ins_486 = regOuts_486;
  assign rport_io_ins_487 = regOuts_487;
  assign rport_io_ins_488 = regOuts_488;
  assign rport_io_ins_489 = regOuts_489;
  assign rport_io_ins_490 = regOuts_490;
  assign rport_io_ins_491 = regOuts_491;
  assign rport_io_ins_492 = regOuts_492;
  assign rport_io_ins_493 = regOuts_493;
  assign rport_io_ins_494 = regOuts_494;
  assign rport_io_ins_495 = regOuts_495;
  assign rport_io_ins_496 = regOuts_496;
  assign rport_io_ins_497 = regOuts_497;
  assign rport_io_ins_498 = regOuts_498;
  assign rport_io_ins_499 = regOuts_499;
  assign rport_io_ins_500 = regOuts_500;
  assign rport_io_ins_501 = regOuts_501;
  assign rport_io_ins_502 = regOuts_502;
  assign rport_io_ins_503 = regOuts_503;
  assign rport_io_ins_504 = regOuts_504;
  assign rport_io_ins_505 = regOuts_505;
  assign rport_io_sel = _T_5611[8:0];
  assign regOuts_0 = regs_0_io_out;
  assign regOuts_1 = regs_1_io_out;
  assign regOuts_2 = regs_2_io_out;
  assign regOuts_3 = regs_3_io_out;
  assign regOuts_4 = regs_4_io_out;
  assign regOuts_5 = regs_5_io_out;
  assign regOuts_6 = regs_6_io_out;
  assign regOuts_7 = regs_7_io_out;
  assign regOuts_8 = regs_8_io_out;
  assign regOuts_9 = regs_9_io_out;
  assign regOuts_10 = regs_10_io_out;
  assign regOuts_11 = regs_11_io_out;
  assign regOuts_12 = regs_12_io_out;
  assign regOuts_13 = regs_13_io_out;
  assign regOuts_14 = regs_14_io_out;
  assign regOuts_15 = regs_15_io_out;
  assign regOuts_16 = regs_16_io_out;
  assign regOuts_17 = regs_17_io_out;
  assign regOuts_18 = regs_18_io_out;
  assign regOuts_19 = regs_19_io_out;
  assign regOuts_20 = regs_20_io_out;
  assign regOuts_21 = regs_21_io_out;
  assign regOuts_22 = regs_22_io_out;
  assign regOuts_23 = regs_23_io_out;
  assign regOuts_24 = regs_24_io_out;
  assign regOuts_25 = regs_25_io_out;
  assign regOuts_26 = regs_26_io_out;
  assign regOuts_27 = regs_27_io_out;
  assign regOuts_28 = regs_28_io_out;
  assign regOuts_29 = regs_29_io_out;
  assign regOuts_30 = regs_30_io_out;
  assign regOuts_31 = regs_31_io_out;
  assign regOuts_32 = regs_32_io_out;
  assign regOuts_33 = regs_33_io_out;
  assign regOuts_34 = regs_34_io_out;
  assign regOuts_35 = regs_35_io_out;
  assign regOuts_36 = regs_36_io_out;
  assign regOuts_37 = regs_37_io_out;
  assign regOuts_38 = regs_38_io_out;
  assign regOuts_39 = regs_39_io_out;
  assign regOuts_40 = regs_40_io_out;
  assign regOuts_41 = regs_41_io_out;
  assign regOuts_42 = regs_42_io_out;
  assign regOuts_43 = regs_43_io_out;
  assign regOuts_44 = regs_44_io_out;
  assign regOuts_45 = regs_45_io_out;
  assign regOuts_46 = regs_46_io_out;
  assign regOuts_47 = regs_47_io_out;
  assign regOuts_48 = regs_48_io_out;
  assign regOuts_49 = regs_49_io_out;
  assign regOuts_50 = regs_50_io_out;
  assign regOuts_51 = regs_51_io_out;
  assign regOuts_52 = regs_52_io_out;
  assign regOuts_53 = regs_53_io_out;
  assign regOuts_54 = regs_54_io_out;
  assign regOuts_55 = regs_55_io_out;
  assign regOuts_56 = regs_56_io_out;
  assign regOuts_57 = regs_57_io_out;
  assign regOuts_58 = regs_58_io_out;
  assign regOuts_59 = regs_59_io_out;
  assign regOuts_60 = regs_60_io_out;
  assign regOuts_61 = regs_61_io_out;
  assign regOuts_62 = regs_62_io_out;
  assign regOuts_63 = regs_63_io_out;
  assign regOuts_64 = regs_64_io_out;
  assign regOuts_65 = regs_65_io_out;
  assign regOuts_66 = regs_66_io_out;
  assign regOuts_67 = regs_67_io_out;
  assign regOuts_68 = regs_68_io_out;
  assign regOuts_69 = regs_69_io_out;
  assign regOuts_70 = regs_70_io_out;
  assign regOuts_71 = regs_71_io_out;
  assign regOuts_72 = regs_72_io_out;
  assign regOuts_73 = regs_73_io_out;
  assign regOuts_74 = regs_74_io_out;
  assign regOuts_75 = regs_75_io_out;
  assign regOuts_76 = regs_76_io_out;
  assign regOuts_77 = regs_77_io_out;
  assign regOuts_78 = regs_78_io_out;
  assign regOuts_79 = regs_79_io_out;
  assign regOuts_80 = regs_80_io_out;
  assign regOuts_81 = regs_81_io_out;
  assign regOuts_82 = regs_82_io_out;
  assign regOuts_83 = regs_83_io_out;
  assign regOuts_84 = regs_84_io_out;
  assign regOuts_85 = regs_85_io_out;
  assign regOuts_86 = regs_86_io_out;
  assign regOuts_87 = regs_87_io_out;
  assign regOuts_88 = regs_88_io_out;
  assign regOuts_89 = regs_89_io_out;
  assign regOuts_90 = regs_90_io_out;
  assign regOuts_91 = regs_91_io_out;
  assign regOuts_92 = regs_92_io_out;
  assign regOuts_93 = regs_93_io_out;
  assign regOuts_94 = regs_94_io_out;
  assign regOuts_95 = regs_95_io_out;
  assign regOuts_96 = regs_96_io_out;
  assign regOuts_97 = regs_97_io_out;
  assign regOuts_98 = regs_98_io_out;
  assign regOuts_99 = regs_99_io_out;
  assign regOuts_100 = regs_100_io_out;
  assign regOuts_101 = regs_101_io_out;
  assign regOuts_102 = regs_102_io_out;
  assign regOuts_103 = regs_103_io_out;
  assign regOuts_104 = regs_104_io_out;
  assign regOuts_105 = regs_105_io_out;
  assign regOuts_106 = regs_106_io_out;
  assign regOuts_107 = regs_107_io_out;
  assign regOuts_108 = regs_108_io_out;
  assign regOuts_109 = regs_109_io_out;
  assign regOuts_110 = regs_110_io_out;
  assign regOuts_111 = regs_111_io_out;
  assign regOuts_112 = regs_112_io_out;
  assign regOuts_113 = regs_113_io_out;
  assign regOuts_114 = regs_114_io_out;
  assign regOuts_115 = regs_115_io_out;
  assign regOuts_116 = regs_116_io_out;
  assign regOuts_117 = regs_117_io_out;
  assign regOuts_118 = regs_118_io_out;
  assign regOuts_119 = regs_119_io_out;
  assign regOuts_120 = regs_120_io_out;
  assign regOuts_121 = regs_121_io_out;
  assign regOuts_122 = regs_122_io_out;
  assign regOuts_123 = regs_123_io_out;
  assign regOuts_124 = regs_124_io_out;
  assign regOuts_125 = regs_125_io_out;
  assign regOuts_126 = regs_126_io_out;
  assign regOuts_127 = regs_127_io_out;
  assign regOuts_128 = regs_128_io_out;
  assign regOuts_129 = regs_129_io_out;
  assign regOuts_130 = regs_130_io_out;
  assign regOuts_131 = regs_131_io_out;
  assign regOuts_132 = regs_132_io_out;
  assign regOuts_133 = regs_133_io_out;
  assign regOuts_134 = regs_134_io_out;
  assign regOuts_135 = regs_135_io_out;
  assign regOuts_136 = regs_136_io_out;
  assign regOuts_137 = regs_137_io_out;
  assign regOuts_138 = regs_138_io_out;
  assign regOuts_139 = regs_139_io_out;
  assign regOuts_140 = regs_140_io_out;
  assign regOuts_141 = regs_141_io_out;
  assign regOuts_142 = regs_142_io_out;
  assign regOuts_143 = regs_143_io_out;
  assign regOuts_144 = regs_144_io_out;
  assign regOuts_145 = regs_145_io_out;
  assign regOuts_146 = regs_146_io_out;
  assign regOuts_147 = regs_147_io_out;
  assign regOuts_148 = regs_148_io_out;
  assign regOuts_149 = regs_149_io_out;
  assign regOuts_150 = regs_150_io_out;
  assign regOuts_151 = regs_151_io_out;
  assign regOuts_152 = regs_152_io_out;
  assign regOuts_153 = regs_153_io_out;
  assign regOuts_154 = regs_154_io_out;
  assign regOuts_155 = regs_155_io_out;
  assign regOuts_156 = regs_156_io_out;
  assign regOuts_157 = regs_157_io_out;
  assign regOuts_158 = regs_158_io_out;
  assign regOuts_159 = regs_159_io_out;
  assign regOuts_160 = regs_160_io_out;
  assign regOuts_161 = regs_161_io_out;
  assign regOuts_162 = regs_162_io_out;
  assign regOuts_163 = regs_163_io_out;
  assign regOuts_164 = regs_164_io_out;
  assign regOuts_165 = regs_165_io_out;
  assign regOuts_166 = regs_166_io_out;
  assign regOuts_167 = regs_167_io_out;
  assign regOuts_168 = regs_168_io_out;
  assign regOuts_169 = regs_169_io_out;
  assign regOuts_170 = regs_170_io_out;
  assign regOuts_171 = regs_171_io_out;
  assign regOuts_172 = regs_172_io_out;
  assign regOuts_173 = regs_173_io_out;
  assign regOuts_174 = regs_174_io_out;
  assign regOuts_175 = regs_175_io_out;
  assign regOuts_176 = regs_176_io_out;
  assign regOuts_177 = regs_177_io_out;
  assign regOuts_178 = regs_178_io_out;
  assign regOuts_179 = regs_179_io_out;
  assign regOuts_180 = regs_180_io_out;
  assign regOuts_181 = regs_181_io_out;
  assign regOuts_182 = regs_182_io_out;
  assign regOuts_183 = regs_183_io_out;
  assign regOuts_184 = regs_184_io_out;
  assign regOuts_185 = regs_185_io_out;
  assign regOuts_186 = regs_186_io_out;
  assign regOuts_187 = regs_187_io_out;
  assign regOuts_188 = regs_188_io_out;
  assign regOuts_189 = regs_189_io_out;
  assign regOuts_190 = regs_190_io_out;
  assign regOuts_191 = regs_191_io_out;
  assign regOuts_192 = regs_192_io_out;
  assign regOuts_193 = regs_193_io_out;
  assign regOuts_194 = regs_194_io_out;
  assign regOuts_195 = regs_195_io_out;
  assign regOuts_196 = regs_196_io_out;
  assign regOuts_197 = regs_197_io_out;
  assign regOuts_198 = regs_198_io_out;
  assign regOuts_199 = regs_199_io_out;
  assign regOuts_200 = regs_200_io_out;
  assign regOuts_201 = regs_201_io_out;
  assign regOuts_202 = regs_202_io_out;
  assign regOuts_203 = regs_203_io_out;
  assign regOuts_204 = regs_204_io_out;
  assign regOuts_205 = regs_205_io_out;
  assign regOuts_206 = regs_206_io_out;
  assign regOuts_207 = regs_207_io_out;
  assign regOuts_208 = regs_208_io_out;
  assign regOuts_209 = regs_209_io_out;
  assign regOuts_210 = regs_210_io_out;
  assign regOuts_211 = regs_211_io_out;
  assign regOuts_212 = regs_212_io_out;
  assign regOuts_213 = regs_213_io_out;
  assign regOuts_214 = regs_214_io_out;
  assign regOuts_215 = regs_215_io_out;
  assign regOuts_216 = regs_216_io_out;
  assign regOuts_217 = regs_217_io_out;
  assign regOuts_218 = regs_218_io_out;
  assign regOuts_219 = regs_219_io_out;
  assign regOuts_220 = regs_220_io_out;
  assign regOuts_221 = regs_221_io_out;
  assign regOuts_222 = regs_222_io_out;
  assign regOuts_223 = regs_223_io_out;
  assign regOuts_224 = regs_224_io_out;
  assign regOuts_225 = regs_225_io_out;
  assign regOuts_226 = regs_226_io_out;
  assign regOuts_227 = regs_227_io_out;
  assign regOuts_228 = regs_228_io_out;
  assign regOuts_229 = regs_229_io_out;
  assign regOuts_230 = regs_230_io_out;
  assign regOuts_231 = regs_231_io_out;
  assign regOuts_232 = regs_232_io_out;
  assign regOuts_233 = regs_233_io_out;
  assign regOuts_234 = regs_234_io_out;
  assign regOuts_235 = regs_235_io_out;
  assign regOuts_236 = regs_236_io_out;
  assign regOuts_237 = regs_237_io_out;
  assign regOuts_238 = regs_238_io_out;
  assign regOuts_239 = regs_239_io_out;
  assign regOuts_240 = regs_240_io_out;
  assign regOuts_241 = regs_241_io_out;
  assign regOuts_242 = regs_242_io_out;
  assign regOuts_243 = regs_243_io_out;
  assign regOuts_244 = regs_244_io_out;
  assign regOuts_245 = regs_245_io_out;
  assign regOuts_246 = regs_246_io_out;
  assign regOuts_247 = regs_247_io_out;
  assign regOuts_248 = regs_248_io_out;
  assign regOuts_249 = regs_249_io_out;
  assign regOuts_250 = regs_250_io_out;
  assign regOuts_251 = regs_251_io_out;
  assign regOuts_252 = regs_252_io_out;
  assign regOuts_253 = regs_253_io_out;
  assign regOuts_254 = regs_254_io_out;
  assign regOuts_255 = regs_255_io_out;
  assign regOuts_256 = regs_256_io_out;
  assign regOuts_257 = regs_257_io_out;
  assign regOuts_258 = regs_258_io_out;
  assign regOuts_259 = regs_259_io_out;
  assign regOuts_260 = regs_260_io_out;
  assign regOuts_261 = regs_261_io_out;
  assign regOuts_262 = regs_262_io_out;
  assign regOuts_263 = regs_263_io_out;
  assign regOuts_264 = regs_264_io_out;
  assign regOuts_265 = regs_265_io_out;
  assign regOuts_266 = regs_266_io_out;
  assign regOuts_267 = regs_267_io_out;
  assign regOuts_268 = regs_268_io_out;
  assign regOuts_269 = regs_269_io_out;
  assign regOuts_270 = regs_270_io_out;
  assign regOuts_271 = regs_271_io_out;
  assign regOuts_272 = regs_272_io_out;
  assign regOuts_273 = regs_273_io_out;
  assign regOuts_274 = regs_274_io_out;
  assign regOuts_275 = regs_275_io_out;
  assign regOuts_276 = regs_276_io_out;
  assign regOuts_277 = regs_277_io_out;
  assign regOuts_278 = regs_278_io_out;
  assign regOuts_279 = regs_279_io_out;
  assign regOuts_280 = regs_280_io_out;
  assign regOuts_281 = regs_281_io_out;
  assign regOuts_282 = regs_282_io_out;
  assign regOuts_283 = regs_283_io_out;
  assign regOuts_284 = regs_284_io_out;
  assign regOuts_285 = regs_285_io_out;
  assign regOuts_286 = regs_286_io_out;
  assign regOuts_287 = regs_287_io_out;
  assign regOuts_288 = regs_288_io_out;
  assign regOuts_289 = regs_289_io_out;
  assign regOuts_290 = regs_290_io_out;
  assign regOuts_291 = regs_291_io_out;
  assign regOuts_292 = regs_292_io_out;
  assign regOuts_293 = regs_293_io_out;
  assign regOuts_294 = regs_294_io_out;
  assign regOuts_295 = regs_295_io_out;
  assign regOuts_296 = regs_296_io_out;
  assign regOuts_297 = regs_297_io_out;
  assign regOuts_298 = regs_298_io_out;
  assign regOuts_299 = regs_299_io_out;
  assign regOuts_300 = regs_300_io_out;
  assign regOuts_301 = regs_301_io_out;
  assign regOuts_302 = regs_302_io_out;
  assign regOuts_303 = regs_303_io_out;
  assign regOuts_304 = regs_304_io_out;
  assign regOuts_305 = regs_305_io_out;
  assign regOuts_306 = regs_306_io_out;
  assign regOuts_307 = regs_307_io_out;
  assign regOuts_308 = regs_308_io_out;
  assign regOuts_309 = regs_309_io_out;
  assign regOuts_310 = regs_310_io_out;
  assign regOuts_311 = regs_311_io_out;
  assign regOuts_312 = regs_312_io_out;
  assign regOuts_313 = regs_313_io_out;
  assign regOuts_314 = regs_314_io_out;
  assign regOuts_315 = regs_315_io_out;
  assign regOuts_316 = regs_316_io_out;
  assign regOuts_317 = regs_317_io_out;
  assign regOuts_318 = regs_318_io_out;
  assign regOuts_319 = regs_319_io_out;
  assign regOuts_320 = regs_320_io_out;
  assign regOuts_321 = regs_321_io_out;
  assign regOuts_322 = regs_322_io_out;
  assign regOuts_323 = regs_323_io_out;
  assign regOuts_324 = regs_324_io_out;
  assign regOuts_325 = regs_325_io_out;
  assign regOuts_326 = regs_326_io_out;
  assign regOuts_327 = regs_327_io_out;
  assign regOuts_328 = regs_328_io_out;
  assign regOuts_329 = regs_329_io_out;
  assign regOuts_330 = regs_330_io_out;
  assign regOuts_331 = regs_331_io_out;
  assign regOuts_332 = regs_332_io_out;
  assign regOuts_333 = regs_333_io_out;
  assign regOuts_334 = regs_334_io_out;
  assign regOuts_335 = regs_335_io_out;
  assign regOuts_336 = regs_336_io_out;
  assign regOuts_337 = regs_337_io_out;
  assign regOuts_338 = regs_338_io_out;
  assign regOuts_339 = regs_339_io_out;
  assign regOuts_340 = regs_340_io_out;
  assign regOuts_341 = regs_341_io_out;
  assign regOuts_342 = regs_342_io_out;
  assign regOuts_343 = regs_343_io_out;
  assign regOuts_344 = regs_344_io_out;
  assign regOuts_345 = regs_345_io_out;
  assign regOuts_346 = regs_346_io_out;
  assign regOuts_347 = regs_347_io_out;
  assign regOuts_348 = regs_348_io_out;
  assign regOuts_349 = regs_349_io_out;
  assign regOuts_350 = regs_350_io_out;
  assign regOuts_351 = regs_351_io_out;
  assign regOuts_352 = regs_352_io_out;
  assign regOuts_353 = regs_353_io_out;
  assign regOuts_354 = regs_354_io_out;
  assign regOuts_355 = regs_355_io_out;
  assign regOuts_356 = regs_356_io_out;
  assign regOuts_357 = regs_357_io_out;
  assign regOuts_358 = regs_358_io_out;
  assign regOuts_359 = regs_359_io_out;
  assign regOuts_360 = regs_360_io_out;
  assign regOuts_361 = regs_361_io_out;
  assign regOuts_362 = regs_362_io_out;
  assign regOuts_363 = regs_363_io_out;
  assign regOuts_364 = regs_364_io_out;
  assign regOuts_365 = regs_365_io_out;
  assign regOuts_366 = regs_366_io_out;
  assign regOuts_367 = regs_367_io_out;
  assign regOuts_368 = regs_368_io_out;
  assign regOuts_369 = regs_369_io_out;
  assign regOuts_370 = regs_370_io_out;
  assign regOuts_371 = regs_371_io_out;
  assign regOuts_372 = regs_372_io_out;
  assign regOuts_373 = regs_373_io_out;
  assign regOuts_374 = regs_374_io_out;
  assign regOuts_375 = regs_375_io_out;
  assign regOuts_376 = regs_376_io_out;
  assign regOuts_377 = regs_377_io_out;
  assign regOuts_378 = regs_378_io_out;
  assign regOuts_379 = regs_379_io_out;
  assign regOuts_380 = regs_380_io_out;
  assign regOuts_381 = regs_381_io_out;
  assign regOuts_382 = regs_382_io_out;
  assign regOuts_383 = regs_383_io_out;
  assign regOuts_384 = regs_384_io_out;
  assign regOuts_385 = regs_385_io_out;
  assign regOuts_386 = regs_386_io_out;
  assign regOuts_387 = regs_387_io_out;
  assign regOuts_388 = regs_388_io_out;
  assign regOuts_389 = regs_389_io_out;
  assign regOuts_390 = regs_390_io_out;
  assign regOuts_391 = regs_391_io_out;
  assign regOuts_392 = regs_392_io_out;
  assign regOuts_393 = regs_393_io_out;
  assign regOuts_394 = regs_394_io_out;
  assign regOuts_395 = regs_395_io_out;
  assign regOuts_396 = regs_396_io_out;
  assign regOuts_397 = regs_397_io_out;
  assign regOuts_398 = regs_398_io_out;
  assign regOuts_399 = regs_399_io_out;
  assign regOuts_400 = regs_400_io_out;
  assign regOuts_401 = regs_401_io_out;
  assign regOuts_402 = regs_402_io_out;
  assign regOuts_403 = regs_403_io_out;
  assign regOuts_404 = regs_404_io_out;
  assign regOuts_405 = regs_405_io_out;
  assign regOuts_406 = regs_406_io_out;
  assign regOuts_407 = regs_407_io_out;
  assign regOuts_408 = regs_408_io_out;
  assign regOuts_409 = regs_409_io_out;
  assign regOuts_410 = regs_410_io_out;
  assign regOuts_411 = regs_411_io_out;
  assign regOuts_412 = regs_412_io_out;
  assign regOuts_413 = regs_413_io_out;
  assign regOuts_414 = regs_414_io_out;
  assign regOuts_415 = regs_415_io_out;
  assign regOuts_416 = regs_416_io_out;
  assign regOuts_417 = regs_417_io_out;
  assign regOuts_418 = regs_418_io_out;
  assign regOuts_419 = regs_419_io_out;
  assign regOuts_420 = regs_420_io_out;
  assign regOuts_421 = regs_421_io_out;
  assign regOuts_422 = regs_422_io_out;
  assign regOuts_423 = regs_423_io_out;
  assign regOuts_424 = regs_424_io_out;
  assign regOuts_425 = regs_425_io_out;
  assign regOuts_426 = regs_426_io_out;
  assign regOuts_427 = regs_427_io_out;
  assign regOuts_428 = regs_428_io_out;
  assign regOuts_429 = regs_429_io_out;
  assign regOuts_430 = regs_430_io_out;
  assign regOuts_431 = regs_431_io_out;
  assign regOuts_432 = regs_432_io_out;
  assign regOuts_433 = regs_433_io_out;
  assign regOuts_434 = regs_434_io_out;
  assign regOuts_435 = regs_435_io_out;
  assign regOuts_436 = regs_436_io_out;
  assign regOuts_437 = regs_437_io_out;
  assign regOuts_438 = regs_438_io_out;
  assign regOuts_439 = regs_439_io_out;
  assign regOuts_440 = regs_440_io_out;
  assign regOuts_441 = regs_441_io_out;
  assign regOuts_442 = regs_442_io_out;
  assign regOuts_443 = regs_443_io_out;
  assign regOuts_444 = regs_444_io_out;
  assign regOuts_445 = regs_445_io_out;
  assign regOuts_446 = regs_446_io_out;
  assign regOuts_447 = regs_447_io_out;
  assign regOuts_448 = regs_448_io_out;
  assign regOuts_449 = regs_449_io_out;
  assign regOuts_450 = regs_450_io_out;
  assign regOuts_451 = regs_451_io_out;
  assign regOuts_452 = regs_452_io_out;
  assign regOuts_453 = regs_453_io_out;
  assign regOuts_454 = regs_454_io_out;
  assign regOuts_455 = regs_455_io_out;
  assign regOuts_456 = regs_456_io_out;
  assign regOuts_457 = regs_457_io_out;
  assign regOuts_458 = regs_458_io_out;
  assign regOuts_459 = regs_459_io_out;
  assign regOuts_460 = regs_460_io_out;
  assign regOuts_461 = regs_461_io_out;
  assign regOuts_462 = regs_462_io_out;
  assign regOuts_463 = regs_463_io_out;
  assign regOuts_464 = regs_464_io_out;
  assign regOuts_465 = regs_465_io_out;
  assign regOuts_466 = regs_466_io_out;
  assign regOuts_467 = regs_467_io_out;
  assign regOuts_468 = regs_468_io_out;
  assign regOuts_469 = regs_469_io_out;
  assign regOuts_470 = regs_470_io_out;
  assign regOuts_471 = regs_471_io_out;
  assign regOuts_472 = regs_472_io_out;
  assign regOuts_473 = regs_473_io_out;
  assign regOuts_474 = regs_474_io_out;
  assign regOuts_475 = regs_475_io_out;
  assign regOuts_476 = regs_476_io_out;
  assign regOuts_477 = regs_477_io_out;
  assign regOuts_478 = regs_478_io_out;
  assign regOuts_479 = regs_479_io_out;
  assign regOuts_480 = regs_480_io_out;
  assign regOuts_481 = regs_481_io_out;
  assign regOuts_482 = regs_482_io_out;
  assign regOuts_483 = regs_483_io_out;
  assign regOuts_484 = regs_484_io_out;
  assign regOuts_485 = regs_485_io_out;
  assign regOuts_486 = regs_486_io_out;
  assign regOuts_487 = regs_487_io_out;
  assign regOuts_488 = regs_488_io_out;
  assign regOuts_489 = regs_489_io_out;
  assign regOuts_490 = regs_490_io_out;
  assign regOuts_491 = regs_491_io_out;
  assign regOuts_492 = regs_492_io_out;
  assign regOuts_493 = regs_493_io_out;
  assign regOuts_494 = regs_494_io_out;
  assign regOuts_495 = regs_495_io_out;
  assign regOuts_496 = regs_496_io_out;
  assign regOuts_497 = regs_497_io_out;
  assign regOuts_498 = regs_498_io_out;
  assign regOuts_499 = regs_499_io_out;
  assign regOuts_500 = regs_500_io_out;
  assign regOuts_501 = regs_501_io_out;
  assign regOuts_502 = regs_502_io_out;
  assign regOuts_503 = regs_503_io_out;
  assign regOuts_504 = regs_504_io_out;
  assign regOuts_505 = regs_505_io_out;
  assign _T_5618_0 = regOuts_0;
  assign _T_5618_1 = regOuts_1;
  assign _T_5618_2 = regOuts_2;
  assign _T_5618_3 = regOuts_3;
  assign _T_5618_4 = regOuts_4;
endmodule
module RetimeWrapper_1798(
  input         clock,
  input         reset,
  input  [39:0] io_in,
  output [39:0] io_out
);
  wire [39:0] sr_out;
  wire [39:0] sr_in;
  wire  sr_flow;
  wire  sr_reset;
  wire  sr_clock;
  RetimeShiftRegister #(.WIDTH(40), .STAGES(1)) sr (
    .out(sr_out),
    .in(sr_in),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out;
  assign sr_in = io_in;
  assign sr_flow = 1'h1;
  assign sr_reset = reset;
  assign sr_clock = clock;
endmodule
module FF_1369(
  input         clock,
  input         reset,
  input  [39:0] io_in,
  output [39:0] io_out,
  input         io_enable
);
  wire [39:0] d;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire [39:0] RetimeWrapper_io_in;
  wire [39:0] RetimeWrapper_io_out;
  wire [39:0] _T_11;
  wire [39:0] _GEN_1;
  RetimeWrapper_1798 RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _GEN_1 = io_enable ? io_in : _T_11;
  assign io_out = _T_11;
  assign d = _GEN_1;
  assign RetimeWrapper_io_in = d;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_11 = RetimeWrapper_io_out;
endmodule
module Counter_443(
  input   clock,
  input   reset,
  input   io_enable,
  output  io_done
);
  wire  reg$_clock;
  wire  reg$_reset;
  wire [39:0] reg$_io_in;
  wire [39:0] reg$_io_out;
  wire  reg$_io_enable;
  wire [40:0] count;
  wire [41:0] _T_13;
  wire [40:0] newval;
  wire  isMax;
  wire [40:0] next;
  wire  _T_15;
  FF_1369 reg$ (
    .clock(reg$_clock),
    .reset(reg$_reset),
    .io_in(reg$_io_in),
    .io_out(reg$_io_out),
    .io_enable(reg$_io_enable)
  );
  assign count = {1'h0,reg$_io_out};
  assign _T_13 = count + 41'h1;
  assign newval = _T_13[40:0];
  assign isMax = newval >= 41'h2cb417800;
  assign next = isMax ? count : newval;
  assign _T_15 = io_enable & isMax;
  assign io_done = _T_15;
  assign reg$_io_in = next[39:0];
  assign reg$_io_enable = io_enable;
  assign reg$_clock = clock;
  assign reg$_reset = reset;
endmodule
module Fringe(
  input          clock,
  input          reset,
  input  [31:0]  io_raddr,
  input          io_wen,
  input  [31:0]  io_waddr,
  input  [63:0]  io_wdata,
  output [63:0]  io_rdata,
  output         io_enable,
  input          io_done,
  output         io_reset,
  output [63:0]  io_argIns_0,
  output [63:0]  io_argIns_1,
  output [63:0]  io_argIns_2,
  input          io_argOuts_0_valid,
  input  [63:0]  io_argOuts_0_bits,
  output         io_memStreams_loads_3_cmd_ready,
  input          io_memStreams_loads_3_cmd_valid,
  input  [63:0]  io_memStreams_loads_3_cmd_bits_addr,
  input          io_memStreams_loads_3_cmd_bits_isWr,
  input  [15:0]  io_memStreams_loads_3_cmd_bits_size,
  input          io_memStreams_loads_3_rdata_ready,
  output         io_memStreams_loads_3_rdata_valid,
  output [31:0]  io_memStreams_loads_3_rdata_bits_0,
  output         io_memStreams_loads_2_cmd_ready,
  input          io_memStreams_loads_2_cmd_valid,
  input  [63:0]  io_memStreams_loads_2_cmd_bits_addr,
  input          io_memStreams_loads_2_cmd_bits_isWr,
  input  [15:0]  io_memStreams_loads_2_cmd_bits_size,
  input          io_memStreams_loads_2_rdata_ready,
  output         io_memStreams_loads_2_rdata_valid,
  output [31:0]  io_memStreams_loads_2_rdata_bits_0,
  output         io_memStreams_loads_1_cmd_ready,
  input          io_memStreams_loads_1_cmd_valid,
  input  [63:0]  io_memStreams_loads_1_cmd_bits_addr,
  input          io_memStreams_loads_1_cmd_bits_isWr,
  input  [15:0]  io_memStreams_loads_1_cmd_bits_size,
  input          io_memStreams_loads_1_rdata_ready,
  output         io_memStreams_loads_1_rdata_valid,
  output [31:0]  io_memStreams_loads_1_rdata_bits_0,
  output         io_memStreams_loads_0_cmd_ready,
  input          io_memStreams_loads_0_cmd_valid,
  input  [63:0]  io_memStreams_loads_0_cmd_bits_addr,
  input          io_memStreams_loads_0_cmd_bits_isWr,
  input  [15:0]  io_memStreams_loads_0_cmd_bits_size,
  input          io_memStreams_loads_0_rdata_ready,
  output         io_memStreams_loads_0_rdata_valid,
  output [31:0]  io_memStreams_loads_0_rdata_bits_0,
  input          io_dram_0_cmd_ready,
  output         io_dram_0_cmd_valid,
  output [63:0]  io_dram_0_cmd_bits_addr,
  output [31:0]  io_dram_0_cmd_bits_size,
  output         io_dram_0_cmd_bits_isWr,
  output [25:0]  io_dram_0_cmd_bits_tag_uid,
  output [5:0]   io_dram_0_cmd_bits_tag_streamId,
  input          io_dram_0_wdata_ready,
  output         io_dram_0_wdata_valid,
  output [31:0]  io_dram_0_wdata_bits_wdata_0,
  output [31:0]  io_dram_0_wdata_bits_wdata_1,
  output [31:0]  io_dram_0_wdata_bits_wdata_2,
  output [31:0]  io_dram_0_wdata_bits_wdata_3,
  output [31:0]  io_dram_0_wdata_bits_wdata_4,
  output [31:0]  io_dram_0_wdata_bits_wdata_5,
  output [31:0]  io_dram_0_wdata_bits_wdata_6,
  output [31:0]  io_dram_0_wdata_bits_wdata_7,
  output [31:0]  io_dram_0_wdata_bits_wdata_8,
  output [31:0]  io_dram_0_wdata_bits_wdata_9,
  output [31:0]  io_dram_0_wdata_bits_wdata_10,
  output [31:0]  io_dram_0_wdata_bits_wdata_11,
  output [31:0]  io_dram_0_wdata_bits_wdata_12,
  output [31:0]  io_dram_0_wdata_bits_wdata_13,
  output [31:0]  io_dram_0_wdata_bits_wdata_14,
  output [31:0]  io_dram_0_wdata_bits_wdata_15,
  output         io_dram_0_wdata_bits_wstrb_0,
  output         io_dram_0_wdata_bits_wstrb_1,
  output         io_dram_0_wdata_bits_wstrb_2,
  output         io_dram_0_wdata_bits_wstrb_3,
  output         io_dram_0_wdata_bits_wstrb_4,
  output         io_dram_0_wdata_bits_wstrb_5,
  output         io_dram_0_wdata_bits_wstrb_6,
  output         io_dram_0_wdata_bits_wstrb_7,
  output         io_dram_0_wdata_bits_wstrb_8,
  output         io_dram_0_wdata_bits_wstrb_9,
  output         io_dram_0_wdata_bits_wstrb_10,
  output         io_dram_0_wdata_bits_wstrb_11,
  output         io_dram_0_wdata_bits_wstrb_12,
  output         io_dram_0_wdata_bits_wstrb_13,
  output         io_dram_0_wdata_bits_wstrb_14,
  output         io_dram_0_wdata_bits_wstrb_15,
  output         io_dram_0_wdata_bits_wstrb_16,
  output         io_dram_0_wdata_bits_wstrb_17,
  output         io_dram_0_wdata_bits_wstrb_18,
  output         io_dram_0_wdata_bits_wstrb_19,
  output         io_dram_0_wdata_bits_wstrb_20,
  output         io_dram_0_wdata_bits_wstrb_21,
  output         io_dram_0_wdata_bits_wstrb_22,
  output         io_dram_0_wdata_bits_wstrb_23,
  output         io_dram_0_wdata_bits_wstrb_24,
  output         io_dram_0_wdata_bits_wstrb_25,
  output         io_dram_0_wdata_bits_wstrb_26,
  output         io_dram_0_wdata_bits_wstrb_27,
  output         io_dram_0_wdata_bits_wstrb_28,
  output         io_dram_0_wdata_bits_wstrb_29,
  output         io_dram_0_wdata_bits_wstrb_30,
  output         io_dram_0_wdata_bits_wstrb_31,
  output         io_dram_0_wdata_bits_wstrb_32,
  output         io_dram_0_wdata_bits_wstrb_33,
  output         io_dram_0_wdata_bits_wstrb_34,
  output         io_dram_0_wdata_bits_wstrb_35,
  output         io_dram_0_wdata_bits_wstrb_36,
  output         io_dram_0_wdata_bits_wstrb_37,
  output         io_dram_0_wdata_bits_wstrb_38,
  output         io_dram_0_wdata_bits_wstrb_39,
  output         io_dram_0_wdata_bits_wstrb_40,
  output         io_dram_0_wdata_bits_wstrb_41,
  output         io_dram_0_wdata_bits_wstrb_42,
  output         io_dram_0_wdata_bits_wstrb_43,
  output         io_dram_0_wdata_bits_wstrb_44,
  output         io_dram_0_wdata_bits_wstrb_45,
  output         io_dram_0_wdata_bits_wstrb_46,
  output         io_dram_0_wdata_bits_wstrb_47,
  output         io_dram_0_wdata_bits_wstrb_48,
  output         io_dram_0_wdata_bits_wstrb_49,
  output         io_dram_0_wdata_bits_wstrb_50,
  output         io_dram_0_wdata_bits_wstrb_51,
  output         io_dram_0_wdata_bits_wstrb_52,
  output         io_dram_0_wdata_bits_wstrb_53,
  output         io_dram_0_wdata_bits_wstrb_54,
  output         io_dram_0_wdata_bits_wstrb_55,
  output         io_dram_0_wdata_bits_wstrb_56,
  output         io_dram_0_wdata_bits_wstrb_57,
  output         io_dram_0_wdata_bits_wstrb_58,
  output         io_dram_0_wdata_bits_wstrb_59,
  output         io_dram_0_wdata_bits_wstrb_60,
  output         io_dram_0_wdata_bits_wstrb_61,
  output         io_dram_0_wdata_bits_wstrb_62,
  output         io_dram_0_wdata_bits_wstrb_63,
  output         io_dram_0_rresp_ready,
  input          io_dram_0_rresp_valid,
  input  [31:0]  io_dram_0_rresp_bits_rdata_0,
  input  [31:0]  io_dram_0_rresp_bits_rdata_1,
  input  [31:0]  io_dram_0_rresp_bits_rdata_2,
  input  [31:0]  io_dram_0_rresp_bits_rdata_3,
  input  [31:0]  io_dram_0_rresp_bits_rdata_4,
  input  [31:0]  io_dram_0_rresp_bits_rdata_5,
  input  [31:0]  io_dram_0_rresp_bits_rdata_6,
  input  [31:0]  io_dram_0_rresp_bits_rdata_7,
  input  [31:0]  io_dram_0_rresp_bits_rdata_8,
  input  [31:0]  io_dram_0_rresp_bits_rdata_9,
  input  [31:0]  io_dram_0_rresp_bits_rdata_10,
  input  [31:0]  io_dram_0_rresp_bits_rdata_11,
  input  [31:0]  io_dram_0_rresp_bits_rdata_12,
  input  [31:0]  io_dram_0_rresp_bits_rdata_13,
  input  [31:0]  io_dram_0_rresp_bits_rdata_14,
  input  [31:0]  io_dram_0_rresp_bits_rdata_15,
  input  [5:0]   io_dram_0_rresp_bits_tag_streamId,
  output         io_dram_0_wresp_ready,
  input          io_dram_0_wresp_valid,
  input  [5:0]   io_dram_0_wresp_bits_tag_streamId,
  input          io_dram_1_cmd_ready,
  output         io_dram_1_cmd_valid,
  output [63:0]  io_dram_1_cmd_bits_addr,
  output [31:0]  io_dram_1_cmd_bits_size,
  output         io_dram_1_cmd_bits_isWr,
  output [25:0]  io_dram_1_cmd_bits_tag_uid,
  output [5:0]   io_dram_1_cmd_bits_tag_streamId,
  input          io_dram_1_wdata_ready,
  output         io_dram_1_wdata_valid,
  output [31:0]  io_dram_1_wdata_bits_wdata_0,
  output [31:0]  io_dram_1_wdata_bits_wdata_1,
  output [31:0]  io_dram_1_wdata_bits_wdata_2,
  output [31:0]  io_dram_1_wdata_bits_wdata_3,
  output [31:0]  io_dram_1_wdata_bits_wdata_4,
  output [31:0]  io_dram_1_wdata_bits_wdata_5,
  output [31:0]  io_dram_1_wdata_bits_wdata_6,
  output [31:0]  io_dram_1_wdata_bits_wdata_7,
  output [31:0]  io_dram_1_wdata_bits_wdata_8,
  output [31:0]  io_dram_1_wdata_bits_wdata_9,
  output [31:0]  io_dram_1_wdata_bits_wdata_10,
  output [31:0]  io_dram_1_wdata_bits_wdata_11,
  output [31:0]  io_dram_1_wdata_bits_wdata_12,
  output [31:0]  io_dram_1_wdata_bits_wdata_13,
  output [31:0]  io_dram_1_wdata_bits_wdata_14,
  output [31:0]  io_dram_1_wdata_bits_wdata_15,
  output         io_dram_1_wdata_bits_wstrb_0,
  output         io_dram_1_wdata_bits_wstrb_1,
  output         io_dram_1_wdata_bits_wstrb_2,
  output         io_dram_1_wdata_bits_wstrb_3,
  output         io_dram_1_wdata_bits_wstrb_4,
  output         io_dram_1_wdata_bits_wstrb_5,
  output         io_dram_1_wdata_bits_wstrb_6,
  output         io_dram_1_wdata_bits_wstrb_7,
  output         io_dram_1_wdata_bits_wstrb_8,
  output         io_dram_1_wdata_bits_wstrb_9,
  output         io_dram_1_wdata_bits_wstrb_10,
  output         io_dram_1_wdata_bits_wstrb_11,
  output         io_dram_1_wdata_bits_wstrb_12,
  output         io_dram_1_wdata_bits_wstrb_13,
  output         io_dram_1_wdata_bits_wstrb_14,
  output         io_dram_1_wdata_bits_wstrb_15,
  output         io_dram_1_wdata_bits_wstrb_16,
  output         io_dram_1_wdata_bits_wstrb_17,
  output         io_dram_1_wdata_bits_wstrb_18,
  output         io_dram_1_wdata_bits_wstrb_19,
  output         io_dram_1_wdata_bits_wstrb_20,
  output         io_dram_1_wdata_bits_wstrb_21,
  output         io_dram_1_wdata_bits_wstrb_22,
  output         io_dram_1_wdata_bits_wstrb_23,
  output         io_dram_1_wdata_bits_wstrb_24,
  output         io_dram_1_wdata_bits_wstrb_25,
  output         io_dram_1_wdata_bits_wstrb_26,
  output         io_dram_1_wdata_bits_wstrb_27,
  output         io_dram_1_wdata_bits_wstrb_28,
  output         io_dram_1_wdata_bits_wstrb_29,
  output         io_dram_1_wdata_bits_wstrb_30,
  output         io_dram_1_wdata_bits_wstrb_31,
  output         io_dram_1_wdata_bits_wstrb_32,
  output         io_dram_1_wdata_bits_wstrb_33,
  output         io_dram_1_wdata_bits_wstrb_34,
  output         io_dram_1_wdata_bits_wstrb_35,
  output         io_dram_1_wdata_bits_wstrb_36,
  output         io_dram_1_wdata_bits_wstrb_37,
  output         io_dram_1_wdata_bits_wstrb_38,
  output         io_dram_1_wdata_bits_wstrb_39,
  output         io_dram_1_wdata_bits_wstrb_40,
  output         io_dram_1_wdata_bits_wstrb_41,
  output         io_dram_1_wdata_bits_wstrb_42,
  output         io_dram_1_wdata_bits_wstrb_43,
  output         io_dram_1_wdata_bits_wstrb_44,
  output         io_dram_1_wdata_bits_wstrb_45,
  output         io_dram_1_wdata_bits_wstrb_46,
  output         io_dram_1_wdata_bits_wstrb_47,
  output         io_dram_1_wdata_bits_wstrb_48,
  output         io_dram_1_wdata_bits_wstrb_49,
  output         io_dram_1_wdata_bits_wstrb_50,
  output         io_dram_1_wdata_bits_wstrb_51,
  output         io_dram_1_wdata_bits_wstrb_52,
  output         io_dram_1_wdata_bits_wstrb_53,
  output         io_dram_1_wdata_bits_wstrb_54,
  output         io_dram_1_wdata_bits_wstrb_55,
  output         io_dram_1_wdata_bits_wstrb_56,
  output         io_dram_1_wdata_bits_wstrb_57,
  output         io_dram_1_wdata_bits_wstrb_58,
  output         io_dram_1_wdata_bits_wstrb_59,
  output         io_dram_1_wdata_bits_wstrb_60,
  output         io_dram_1_wdata_bits_wstrb_61,
  output         io_dram_1_wdata_bits_wstrb_62,
  output         io_dram_1_wdata_bits_wstrb_63,
  output         io_dram_1_rresp_ready,
  input          io_dram_1_rresp_valid,
  input  [31:0]  io_dram_1_rresp_bits_rdata_0,
  input  [31:0]  io_dram_1_rresp_bits_rdata_1,
  input  [31:0]  io_dram_1_rresp_bits_rdata_2,
  input  [31:0]  io_dram_1_rresp_bits_rdata_3,
  input  [31:0]  io_dram_1_rresp_bits_rdata_4,
  input  [31:0]  io_dram_1_rresp_bits_rdata_5,
  input  [31:0]  io_dram_1_rresp_bits_rdata_6,
  input  [31:0]  io_dram_1_rresp_bits_rdata_7,
  input  [31:0]  io_dram_1_rresp_bits_rdata_8,
  input  [31:0]  io_dram_1_rresp_bits_rdata_9,
  input  [31:0]  io_dram_1_rresp_bits_rdata_10,
  input  [31:0]  io_dram_1_rresp_bits_rdata_11,
  input  [31:0]  io_dram_1_rresp_bits_rdata_12,
  input  [31:0]  io_dram_1_rresp_bits_rdata_13,
  input  [31:0]  io_dram_1_rresp_bits_rdata_14,
  input  [31:0]  io_dram_1_rresp_bits_rdata_15,
  input  [5:0]   io_dram_1_rresp_bits_tag_streamId,
  output         io_dram_1_wresp_ready,
  input          io_dram_1_wresp_valid,
  input  [5:0]   io_dram_1_wresp_bits_tag_streamId,
  input          io_dram_2_cmd_ready,
  output         io_dram_2_cmd_valid,
  output [63:0]  io_dram_2_cmd_bits_addr,
  output [31:0]  io_dram_2_cmd_bits_size,
  output         io_dram_2_cmd_bits_isWr,
  output [25:0]  io_dram_2_cmd_bits_tag_uid,
  output [5:0]   io_dram_2_cmd_bits_tag_streamId,
  input          io_dram_2_wdata_ready,
  output         io_dram_2_wdata_valid,
  output [31:0]  io_dram_2_wdata_bits_wdata_0,
  output [31:0]  io_dram_2_wdata_bits_wdata_1,
  output [31:0]  io_dram_2_wdata_bits_wdata_2,
  output [31:0]  io_dram_2_wdata_bits_wdata_3,
  output [31:0]  io_dram_2_wdata_bits_wdata_4,
  output [31:0]  io_dram_2_wdata_bits_wdata_5,
  output [31:0]  io_dram_2_wdata_bits_wdata_6,
  output [31:0]  io_dram_2_wdata_bits_wdata_7,
  output [31:0]  io_dram_2_wdata_bits_wdata_8,
  output [31:0]  io_dram_2_wdata_bits_wdata_9,
  output [31:0]  io_dram_2_wdata_bits_wdata_10,
  output [31:0]  io_dram_2_wdata_bits_wdata_11,
  output [31:0]  io_dram_2_wdata_bits_wdata_12,
  output [31:0]  io_dram_2_wdata_bits_wdata_13,
  output [31:0]  io_dram_2_wdata_bits_wdata_14,
  output [31:0]  io_dram_2_wdata_bits_wdata_15,
  output         io_dram_2_wdata_bits_wstrb_0,
  output         io_dram_2_wdata_bits_wstrb_1,
  output         io_dram_2_wdata_bits_wstrb_2,
  output         io_dram_2_wdata_bits_wstrb_3,
  output         io_dram_2_wdata_bits_wstrb_4,
  output         io_dram_2_wdata_bits_wstrb_5,
  output         io_dram_2_wdata_bits_wstrb_6,
  output         io_dram_2_wdata_bits_wstrb_7,
  output         io_dram_2_wdata_bits_wstrb_8,
  output         io_dram_2_wdata_bits_wstrb_9,
  output         io_dram_2_wdata_bits_wstrb_10,
  output         io_dram_2_wdata_bits_wstrb_11,
  output         io_dram_2_wdata_bits_wstrb_12,
  output         io_dram_2_wdata_bits_wstrb_13,
  output         io_dram_2_wdata_bits_wstrb_14,
  output         io_dram_2_wdata_bits_wstrb_15,
  output         io_dram_2_wdata_bits_wstrb_16,
  output         io_dram_2_wdata_bits_wstrb_17,
  output         io_dram_2_wdata_bits_wstrb_18,
  output         io_dram_2_wdata_bits_wstrb_19,
  output         io_dram_2_wdata_bits_wstrb_20,
  output         io_dram_2_wdata_bits_wstrb_21,
  output         io_dram_2_wdata_bits_wstrb_22,
  output         io_dram_2_wdata_bits_wstrb_23,
  output         io_dram_2_wdata_bits_wstrb_24,
  output         io_dram_2_wdata_bits_wstrb_25,
  output         io_dram_2_wdata_bits_wstrb_26,
  output         io_dram_2_wdata_bits_wstrb_27,
  output         io_dram_2_wdata_bits_wstrb_28,
  output         io_dram_2_wdata_bits_wstrb_29,
  output         io_dram_2_wdata_bits_wstrb_30,
  output         io_dram_2_wdata_bits_wstrb_31,
  output         io_dram_2_wdata_bits_wstrb_32,
  output         io_dram_2_wdata_bits_wstrb_33,
  output         io_dram_2_wdata_bits_wstrb_34,
  output         io_dram_2_wdata_bits_wstrb_35,
  output         io_dram_2_wdata_bits_wstrb_36,
  output         io_dram_2_wdata_bits_wstrb_37,
  output         io_dram_2_wdata_bits_wstrb_38,
  output         io_dram_2_wdata_bits_wstrb_39,
  output         io_dram_2_wdata_bits_wstrb_40,
  output         io_dram_2_wdata_bits_wstrb_41,
  output         io_dram_2_wdata_bits_wstrb_42,
  output         io_dram_2_wdata_bits_wstrb_43,
  output         io_dram_2_wdata_bits_wstrb_44,
  output         io_dram_2_wdata_bits_wstrb_45,
  output         io_dram_2_wdata_bits_wstrb_46,
  output         io_dram_2_wdata_bits_wstrb_47,
  output         io_dram_2_wdata_bits_wstrb_48,
  output         io_dram_2_wdata_bits_wstrb_49,
  output         io_dram_2_wdata_bits_wstrb_50,
  output         io_dram_2_wdata_bits_wstrb_51,
  output         io_dram_2_wdata_bits_wstrb_52,
  output         io_dram_2_wdata_bits_wstrb_53,
  output         io_dram_2_wdata_bits_wstrb_54,
  output         io_dram_2_wdata_bits_wstrb_55,
  output         io_dram_2_wdata_bits_wstrb_56,
  output         io_dram_2_wdata_bits_wstrb_57,
  output         io_dram_2_wdata_bits_wstrb_58,
  output         io_dram_2_wdata_bits_wstrb_59,
  output         io_dram_2_wdata_bits_wstrb_60,
  output         io_dram_2_wdata_bits_wstrb_61,
  output         io_dram_2_wdata_bits_wstrb_62,
  output         io_dram_2_wdata_bits_wstrb_63,
  output         io_dram_2_rresp_ready,
  input          io_dram_2_rresp_valid,
  input  [31:0]  io_dram_2_rresp_bits_rdata_0,
  input  [31:0]  io_dram_2_rresp_bits_rdata_1,
  input  [31:0]  io_dram_2_rresp_bits_rdata_2,
  input  [31:0]  io_dram_2_rresp_bits_rdata_3,
  input  [31:0]  io_dram_2_rresp_bits_rdata_4,
  input  [31:0]  io_dram_2_rresp_bits_rdata_5,
  input  [31:0]  io_dram_2_rresp_bits_rdata_6,
  input  [31:0]  io_dram_2_rresp_bits_rdata_7,
  input  [31:0]  io_dram_2_rresp_bits_rdata_8,
  input  [31:0]  io_dram_2_rresp_bits_rdata_9,
  input  [31:0]  io_dram_2_rresp_bits_rdata_10,
  input  [31:0]  io_dram_2_rresp_bits_rdata_11,
  input  [31:0]  io_dram_2_rresp_bits_rdata_12,
  input  [31:0]  io_dram_2_rresp_bits_rdata_13,
  input  [31:0]  io_dram_2_rresp_bits_rdata_14,
  input  [31:0]  io_dram_2_rresp_bits_rdata_15,
  input  [5:0]   io_dram_2_rresp_bits_tag_streamId,
  output         io_dram_2_wresp_ready,
  input          io_dram_2_wresp_valid,
  input  [5:0]   io_dram_2_wresp_bits_tag_streamId,
  input          io_dram_3_cmd_ready,
  output         io_dram_3_cmd_valid,
  output [63:0]  io_dram_3_cmd_bits_addr,
  output [31:0]  io_dram_3_cmd_bits_size,
  output         io_dram_3_cmd_bits_isWr,
  output [25:0]  io_dram_3_cmd_bits_tag_uid,
  output [5:0]   io_dram_3_cmd_bits_tag_streamId,
  input          io_dram_3_wdata_ready,
  output         io_dram_3_wdata_valid,
  output [31:0]  io_dram_3_wdata_bits_wdata_0,
  output [31:0]  io_dram_3_wdata_bits_wdata_1,
  output [31:0]  io_dram_3_wdata_bits_wdata_2,
  output [31:0]  io_dram_3_wdata_bits_wdata_3,
  output [31:0]  io_dram_3_wdata_bits_wdata_4,
  output [31:0]  io_dram_3_wdata_bits_wdata_5,
  output [31:0]  io_dram_3_wdata_bits_wdata_6,
  output [31:0]  io_dram_3_wdata_bits_wdata_7,
  output [31:0]  io_dram_3_wdata_bits_wdata_8,
  output [31:0]  io_dram_3_wdata_bits_wdata_9,
  output [31:0]  io_dram_3_wdata_bits_wdata_10,
  output [31:0]  io_dram_3_wdata_bits_wdata_11,
  output [31:0]  io_dram_3_wdata_bits_wdata_12,
  output [31:0]  io_dram_3_wdata_bits_wdata_13,
  output [31:0]  io_dram_3_wdata_bits_wdata_14,
  output [31:0]  io_dram_3_wdata_bits_wdata_15,
  output         io_dram_3_wdata_bits_wstrb_0,
  output         io_dram_3_wdata_bits_wstrb_1,
  output         io_dram_3_wdata_bits_wstrb_2,
  output         io_dram_3_wdata_bits_wstrb_3,
  output         io_dram_3_wdata_bits_wstrb_4,
  output         io_dram_3_wdata_bits_wstrb_5,
  output         io_dram_3_wdata_bits_wstrb_6,
  output         io_dram_3_wdata_bits_wstrb_7,
  output         io_dram_3_wdata_bits_wstrb_8,
  output         io_dram_3_wdata_bits_wstrb_9,
  output         io_dram_3_wdata_bits_wstrb_10,
  output         io_dram_3_wdata_bits_wstrb_11,
  output         io_dram_3_wdata_bits_wstrb_12,
  output         io_dram_3_wdata_bits_wstrb_13,
  output         io_dram_3_wdata_bits_wstrb_14,
  output         io_dram_3_wdata_bits_wstrb_15,
  output         io_dram_3_wdata_bits_wstrb_16,
  output         io_dram_3_wdata_bits_wstrb_17,
  output         io_dram_3_wdata_bits_wstrb_18,
  output         io_dram_3_wdata_bits_wstrb_19,
  output         io_dram_3_wdata_bits_wstrb_20,
  output         io_dram_3_wdata_bits_wstrb_21,
  output         io_dram_3_wdata_bits_wstrb_22,
  output         io_dram_3_wdata_bits_wstrb_23,
  output         io_dram_3_wdata_bits_wstrb_24,
  output         io_dram_3_wdata_bits_wstrb_25,
  output         io_dram_3_wdata_bits_wstrb_26,
  output         io_dram_3_wdata_bits_wstrb_27,
  output         io_dram_3_wdata_bits_wstrb_28,
  output         io_dram_3_wdata_bits_wstrb_29,
  output         io_dram_3_wdata_bits_wstrb_30,
  output         io_dram_3_wdata_bits_wstrb_31,
  output         io_dram_3_wdata_bits_wstrb_32,
  output         io_dram_3_wdata_bits_wstrb_33,
  output         io_dram_3_wdata_bits_wstrb_34,
  output         io_dram_3_wdata_bits_wstrb_35,
  output         io_dram_3_wdata_bits_wstrb_36,
  output         io_dram_3_wdata_bits_wstrb_37,
  output         io_dram_3_wdata_bits_wstrb_38,
  output         io_dram_3_wdata_bits_wstrb_39,
  output         io_dram_3_wdata_bits_wstrb_40,
  output         io_dram_3_wdata_bits_wstrb_41,
  output         io_dram_3_wdata_bits_wstrb_42,
  output         io_dram_3_wdata_bits_wstrb_43,
  output         io_dram_3_wdata_bits_wstrb_44,
  output         io_dram_3_wdata_bits_wstrb_45,
  output         io_dram_3_wdata_bits_wstrb_46,
  output         io_dram_3_wdata_bits_wstrb_47,
  output         io_dram_3_wdata_bits_wstrb_48,
  output         io_dram_3_wdata_bits_wstrb_49,
  output         io_dram_3_wdata_bits_wstrb_50,
  output         io_dram_3_wdata_bits_wstrb_51,
  output         io_dram_3_wdata_bits_wstrb_52,
  output         io_dram_3_wdata_bits_wstrb_53,
  output         io_dram_3_wdata_bits_wstrb_54,
  output         io_dram_3_wdata_bits_wstrb_55,
  output         io_dram_3_wdata_bits_wstrb_56,
  output         io_dram_3_wdata_bits_wstrb_57,
  output         io_dram_3_wdata_bits_wstrb_58,
  output         io_dram_3_wdata_bits_wstrb_59,
  output         io_dram_3_wdata_bits_wstrb_60,
  output         io_dram_3_wdata_bits_wstrb_61,
  output         io_dram_3_wdata_bits_wstrb_62,
  output         io_dram_3_wdata_bits_wstrb_63,
  output         io_dram_3_rresp_ready,
  input          io_dram_3_rresp_valid,
  input  [31:0]  io_dram_3_rresp_bits_rdata_0,
  input  [31:0]  io_dram_3_rresp_bits_rdata_1,
  input  [31:0]  io_dram_3_rresp_bits_rdata_2,
  input  [31:0]  io_dram_3_rresp_bits_rdata_3,
  input  [31:0]  io_dram_3_rresp_bits_rdata_4,
  input  [31:0]  io_dram_3_rresp_bits_rdata_5,
  input  [31:0]  io_dram_3_rresp_bits_rdata_6,
  input  [31:0]  io_dram_3_rresp_bits_rdata_7,
  input  [31:0]  io_dram_3_rresp_bits_rdata_8,
  input  [31:0]  io_dram_3_rresp_bits_rdata_9,
  input  [31:0]  io_dram_3_rresp_bits_rdata_10,
  input  [31:0]  io_dram_3_rresp_bits_rdata_11,
  input  [31:0]  io_dram_3_rresp_bits_rdata_12,
  input  [31:0]  io_dram_3_rresp_bits_rdata_13,
  input  [31:0]  io_dram_3_rresp_bits_rdata_14,
  input  [31:0]  io_dram_3_rresp_bits_rdata_15,
  input  [5:0]   io_dram_3_rresp_bits_tag_streamId,
  output         io_dram_3_wresp_ready,
  input          io_dram_3_wresp_valid,
  input  [5:0]   io_dram_3_wresp_bits_tag_streamId,
  input  [63:0]  io_TOP_AXI_AWADDR,
  input  [7:0]   io_TOP_AXI_AWLEN,
  input          io_TOP_AXI_AWVALID,
  input          io_TOP_AXI_AWREADY,
  input          io_TOP_AXI_ARID,
  input  [63:0]  io_TOP_AXI_ARADDR,
  input  [7:0]   io_TOP_AXI_ARLEN,
  input  [2:0]   io_TOP_AXI_ARSIZE,
  input  [1:0]   io_TOP_AXI_ARBURST,
  input          io_TOP_AXI_ARVALID,
  input          io_TOP_AXI_ARREADY,
  input  [511:0] io_TOP_AXI_WDATA,
  input  [63:0]  io_TOP_AXI_WSTRB,
  input          io_TOP_AXI_WVALID,
  input          io_TOP_AXI_WREADY,
  input          io_TOP_AXI_RVALID,
  input          io_TOP_AXI_RREADY,
  input          io_TOP_AXI_BVALID,
  input          io_TOP_AXI_BREADY,
  input  [63:0]  io_DWIDTH_AXI_AWADDR,
  input  [7:0]   io_DWIDTH_AXI_AWLEN,
  input          io_DWIDTH_AXI_AWVALID,
  input          io_DWIDTH_AXI_AWREADY,
  input  [63:0]  io_DWIDTH_AXI_ARADDR,
  input  [7:0]   io_DWIDTH_AXI_ARLEN,
  input  [2:0]   io_DWIDTH_AXI_ARSIZE,
  input  [1:0]   io_DWIDTH_AXI_ARBURST,
  input          io_DWIDTH_AXI_ARVALID,
  input          io_DWIDTH_AXI_ARREADY,
  input  [511:0] io_DWIDTH_AXI_WDATA,
  input  [63:0]  io_DWIDTH_AXI_WSTRB,
  input          io_DWIDTH_AXI_WVALID,
  input          io_DWIDTH_AXI_WREADY,
  input          io_DWIDTH_AXI_RVALID,
  input          io_DWIDTH_AXI_RREADY,
  input          io_DWIDTH_AXI_BVALID,
  input          io_DWIDTH_AXI_BREADY
);
  wire  mags_0_clock;
  wire  mags_0_reset;
  wire  mags_0_io_enable;
  wire  mags_0_io_reset;
  wire  mags_0_io_app_loads_0_cmd_ready;
  wire  mags_0_io_app_loads_0_cmd_valid;
  wire [63:0] mags_0_io_app_loads_0_cmd_bits_addr;
  wire  mags_0_io_app_loads_0_cmd_bits_isWr;
  wire [15:0] mags_0_io_app_loads_0_cmd_bits_size;
  wire  mags_0_io_app_loads_0_rdata_ready;
  wire  mags_0_io_app_loads_0_rdata_valid;
  wire [31:0] mags_0_io_app_loads_0_rdata_bits_0;
  wire  mags_0_io_dram_cmd_ready;
  wire  mags_0_io_dram_cmd_valid;
  wire [63:0] mags_0_io_dram_cmd_bits_addr;
  wire [31:0] mags_0_io_dram_cmd_bits_size;
  wire  mags_0_io_dram_cmd_bits_isWr;
  wire [25:0] mags_0_io_dram_cmd_bits_tag_uid;
  wire [5:0] mags_0_io_dram_cmd_bits_tag_streamId;
  wire  mags_0_io_dram_wdata_ready;
  wire  mags_0_io_dram_wdata_valid;
  wire [31:0] mags_0_io_dram_wdata_bits_wdata_0;
  wire [31:0] mags_0_io_dram_wdata_bits_wdata_1;
  wire [31:0] mags_0_io_dram_wdata_bits_wdata_2;
  wire [31:0] mags_0_io_dram_wdata_bits_wdata_3;
  wire [31:0] mags_0_io_dram_wdata_bits_wdata_4;
  wire [31:0] mags_0_io_dram_wdata_bits_wdata_5;
  wire [31:0] mags_0_io_dram_wdata_bits_wdata_6;
  wire [31:0] mags_0_io_dram_wdata_bits_wdata_7;
  wire [31:0] mags_0_io_dram_wdata_bits_wdata_8;
  wire [31:0] mags_0_io_dram_wdata_bits_wdata_9;
  wire [31:0] mags_0_io_dram_wdata_bits_wdata_10;
  wire [31:0] mags_0_io_dram_wdata_bits_wdata_11;
  wire [31:0] mags_0_io_dram_wdata_bits_wdata_12;
  wire [31:0] mags_0_io_dram_wdata_bits_wdata_13;
  wire [31:0] mags_0_io_dram_wdata_bits_wdata_14;
  wire [31:0] mags_0_io_dram_wdata_bits_wdata_15;
  wire  mags_0_io_dram_wdata_bits_wstrb_0;
  wire  mags_0_io_dram_wdata_bits_wstrb_1;
  wire  mags_0_io_dram_wdata_bits_wstrb_2;
  wire  mags_0_io_dram_wdata_bits_wstrb_3;
  wire  mags_0_io_dram_wdata_bits_wstrb_4;
  wire  mags_0_io_dram_wdata_bits_wstrb_5;
  wire  mags_0_io_dram_wdata_bits_wstrb_6;
  wire  mags_0_io_dram_wdata_bits_wstrb_7;
  wire  mags_0_io_dram_wdata_bits_wstrb_8;
  wire  mags_0_io_dram_wdata_bits_wstrb_9;
  wire  mags_0_io_dram_wdata_bits_wstrb_10;
  wire  mags_0_io_dram_wdata_bits_wstrb_11;
  wire  mags_0_io_dram_wdata_bits_wstrb_12;
  wire  mags_0_io_dram_wdata_bits_wstrb_13;
  wire  mags_0_io_dram_wdata_bits_wstrb_14;
  wire  mags_0_io_dram_wdata_bits_wstrb_15;
  wire  mags_0_io_dram_wdata_bits_wstrb_16;
  wire  mags_0_io_dram_wdata_bits_wstrb_17;
  wire  mags_0_io_dram_wdata_bits_wstrb_18;
  wire  mags_0_io_dram_wdata_bits_wstrb_19;
  wire  mags_0_io_dram_wdata_bits_wstrb_20;
  wire  mags_0_io_dram_wdata_bits_wstrb_21;
  wire  mags_0_io_dram_wdata_bits_wstrb_22;
  wire  mags_0_io_dram_wdata_bits_wstrb_23;
  wire  mags_0_io_dram_wdata_bits_wstrb_24;
  wire  mags_0_io_dram_wdata_bits_wstrb_25;
  wire  mags_0_io_dram_wdata_bits_wstrb_26;
  wire  mags_0_io_dram_wdata_bits_wstrb_27;
  wire  mags_0_io_dram_wdata_bits_wstrb_28;
  wire  mags_0_io_dram_wdata_bits_wstrb_29;
  wire  mags_0_io_dram_wdata_bits_wstrb_30;
  wire  mags_0_io_dram_wdata_bits_wstrb_31;
  wire  mags_0_io_dram_wdata_bits_wstrb_32;
  wire  mags_0_io_dram_wdata_bits_wstrb_33;
  wire  mags_0_io_dram_wdata_bits_wstrb_34;
  wire  mags_0_io_dram_wdata_bits_wstrb_35;
  wire  mags_0_io_dram_wdata_bits_wstrb_36;
  wire  mags_0_io_dram_wdata_bits_wstrb_37;
  wire  mags_0_io_dram_wdata_bits_wstrb_38;
  wire  mags_0_io_dram_wdata_bits_wstrb_39;
  wire  mags_0_io_dram_wdata_bits_wstrb_40;
  wire  mags_0_io_dram_wdata_bits_wstrb_41;
  wire  mags_0_io_dram_wdata_bits_wstrb_42;
  wire  mags_0_io_dram_wdata_bits_wstrb_43;
  wire  mags_0_io_dram_wdata_bits_wstrb_44;
  wire  mags_0_io_dram_wdata_bits_wstrb_45;
  wire  mags_0_io_dram_wdata_bits_wstrb_46;
  wire  mags_0_io_dram_wdata_bits_wstrb_47;
  wire  mags_0_io_dram_wdata_bits_wstrb_48;
  wire  mags_0_io_dram_wdata_bits_wstrb_49;
  wire  mags_0_io_dram_wdata_bits_wstrb_50;
  wire  mags_0_io_dram_wdata_bits_wstrb_51;
  wire  mags_0_io_dram_wdata_bits_wstrb_52;
  wire  mags_0_io_dram_wdata_bits_wstrb_53;
  wire  mags_0_io_dram_wdata_bits_wstrb_54;
  wire  mags_0_io_dram_wdata_bits_wstrb_55;
  wire  mags_0_io_dram_wdata_bits_wstrb_56;
  wire  mags_0_io_dram_wdata_bits_wstrb_57;
  wire  mags_0_io_dram_wdata_bits_wstrb_58;
  wire  mags_0_io_dram_wdata_bits_wstrb_59;
  wire  mags_0_io_dram_wdata_bits_wstrb_60;
  wire  mags_0_io_dram_wdata_bits_wstrb_61;
  wire  mags_0_io_dram_wdata_bits_wstrb_62;
  wire  mags_0_io_dram_wdata_bits_wstrb_63;
  wire  mags_0_io_dram_rresp_ready;
  wire  mags_0_io_dram_rresp_valid;
  wire [31:0] mags_0_io_dram_rresp_bits_rdata_0;
  wire [31:0] mags_0_io_dram_rresp_bits_rdata_1;
  wire [31:0] mags_0_io_dram_rresp_bits_rdata_2;
  wire [31:0] mags_0_io_dram_rresp_bits_rdata_3;
  wire [31:0] mags_0_io_dram_rresp_bits_rdata_4;
  wire [31:0] mags_0_io_dram_rresp_bits_rdata_5;
  wire [31:0] mags_0_io_dram_rresp_bits_rdata_6;
  wire [31:0] mags_0_io_dram_rresp_bits_rdata_7;
  wire [31:0] mags_0_io_dram_rresp_bits_rdata_8;
  wire [31:0] mags_0_io_dram_rresp_bits_rdata_9;
  wire [31:0] mags_0_io_dram_rresp_bits_rdata_10;
  wire [31:0] mags_0_io_dram_rresp_bits_rdata_11;
  wire [31:0] mags_0_io_dram_rresp_bits_rdata_12;
  wire [31:0] mags_0_io_dram_rresp_bits_rdata_13;
  wire [31:0] mags_0_io_dram_rresp_bits_rdata_14;
  wire [31:0] mags_0_io_dram_rresp_bits_rdata_15;
  wire [5:0] mags_0_io_dram_rresp_bits_tag_streamId;
  wire  mags_0_io_dram_wresp_ready;
  wire  mags_0_io_dram_wresp_valid;
  wire [5:0] mags_0_io_dram_wresp_bits_tag_streamId;
  wire [31:0] mags_0_io_debugSignals_0;
  wire [31:0] mags_0_io_debugSignals_1;
  wire [31:0] mags_0_io_debugSignals_2;
  wire [31:0] mags_0_io_debugSignals_3;
  wire [31:0] mags_0_io_debugSignals_4;
  wire [31:0] mags_0_io_debugSignals_5;
  wire [31:0] mags_0_io_debugSignals_6;
  wire [31:0] mags_0_io_debugSignals_7;
  wire [31:0] mags_0_io_debugSignals_8;
  wire [31:0] mags_0_io_debugSignals_9;
  wire [31:0] mags_0_io_debugSignals_10;
  wire [31:0] mags_0_io_debugSignals_11;
  wire [31:0] mags_0_io_debugSignals_12;
  wire [31:0] mags_0_io_debugSignals_13;
  wire [31:0] mags_0_io_debugSignals_14;
  wire [31:0] mags_0_io_debugSignals_15;
  wire [31:0] mags_0_io_debugSignals_16;
  wire [31:0] mags_0_io_debugSignals_17;
  wire [31:0] mags_0_io_debugSignals_18;
  wire [31:0] mags_0_io_debugSignals_19;
  wire [31:0] mags_0_io_debugSignals_20;
  wire [31:0] mags_0_io_debugSignals_21;
  wire [31:0] mags_0_io_debugSignals_22;
  wire [31:0] mags_0_io_debugSignals_23;
  wire [31:0] mags_0_io_debugSignals_24;
  wire [31:0] mags_0_io_debugSignals_25;
  wire [31:0] mags_0_io_debugSignals_26;
  wire [31:0] mags_0_io_debugSignals_27;
  wire [31:0] mags_0_io_debugSignals_28;
  wire [31:0] mags_0_io_debugSignals_29;
  wire [31:0] mags_0_io_debugSignals_30;
  wire [31:0] mags_0_io_debugSignals_31;
  wire [31:0] mags_0_io_debugSignals_32;
  wire [31:0] mags_0_io_debugSignals_33;
  wire [31:0] mags_0_io_debugSignals_34;
  wire [31:0] mags_0_io_debugSignals_35;
  wire [31:0] mags_0_io_debugSignals_36;
  wire [31:0] mags_0_io_debugSignals_37;
  wire [31:0] mags_0_io_debugSignals_38;
  wire [31:0] mags_0_io_debugSignals_39;
  wire [31:0] mags_0_io_debugSignals_40;
  wire [31:0] mags_0_io_debugSignals_41;
  wire [31:0] mags_0_io_debugSignals_42;
  wire [31:0] mags_0_io_debugSignals_43;
  wire [31:0] mags_0_io_debugSignals_44;
  wire [31:0] mags_0_io_debugSignals_45;
  wire [31:0] mags_0_io_debugSignals_46;
  wire [31:0] mags_0_io_debugSignals_47;
  wire [31:0] mags_0_io_debugSignals_48;
  wire [31:0] mags_0_io_debugSignals_49;
  wire [31:0] mags_0_io_debugSignals_50;
  wire [31:0] mags_0_io_debugSignals_51;
  wire [31:0] mags_0_io_debugSignals_52;
  wire [31:0] mags_0_io_debugSignals_53;
  wire [31:0] mags_0_io_debugSignals_54;
  wire [31:0] mags_0_io_debugSignals_55;
  wire [31:0] mags_0_io_debugSignals_56;
  wire [31:0] mags_0_io_debugSignals_57;
  wire [31:0] mags_0_io_debugSignals_58;
  wire [31:0] mags_0_io_debugSignals_59;
  wire [31:0] mags_0_io_debugSignals_60;
  wire [31:0] mags_0_io_debugSignals_61;
  wire [31:0] mags_0_io_debugSignals_62;
  wire [31:0] mags_0_io_debugSignals_63;
  wire [31:0] mags_0_io_debugSignals_64;
  wire [31:0] mags_0_io_debugSignals_65;
  wire [31:0] mags_0_io_debugSignals_66;
  wire [31:0] mags_0_io_debugSignals_67;
  wire [31:0] mags_0_io_debugSignals_68;
  wire [31:0] mags_0_io_debugSignals_69;
  wire [31:0] mags_0_io_debugSignals_70;
  wire [31:0] mags_0_io_debugSignals_71;
  wire [31:0] mags_0_io_debugSignals_72;
  wire [31:0] mags_0_io_debugSignals_73;
  wire [31:0] mags_0_io_debugSignals_74;
  wire [31:0] mags_0_io_debugSignals_75;
  wire [31:0] mags_0_io_debugSignals_76;
  wire [31:0] mags_0_io_debugSignals_77;
  wire [31:0] mags_0_io_debugSignals_78;
  wire [31:0] mags_0_io_debugSignals_79;
  wire [31:0] mags_0_io_debugSignals_80;
  wire [31:0] mags_0_io_debugSignals_81;
  wire [31:0] mags_0_io_debugSignals_82;
  wire [31:0] mags_0_io_debugSignals_83;
  wire [31:0] mags_0_io_debugSignals_84;
  wire [31:0] mags_0_io_debugSignals_85;
  wire [31:0] mags_0_io_debugSignals_86;
  wire [31:0] mags_0_io_debugSignals_87;
  wire [31:0] mags_0_io_debugSignals_88;
  wire [31:0] mags_0_io_debugSignals_89;
  wire [31:0] mags_0_io_debugSignals_90;
  wire [31:0] mags_0_io_debugSignals_91;
  wire [31:0] mags_0_io_debugSignals_92;
  wire [31:0] mags_0_io_debugSignals_93;
  wire [31:0] mags_0_io_debugSignals_94;
  wire [31:0] mags_0_io_debugSignals_95;
  wire [31:0] mags_0_io_debugSignals_96;
  wire [31:0] mags_0_io_debugSignals_97;
  wire [31:0] mags_0_io_debugSignals_98;
  wire [31:0] mags_0_io_debugSignals_99;
  wire [31:0] mags_0_io_debugSignals_100;
  wire [31:0] mags_0_io_debugSignals_101;
  wire [31:0] mags_0_io_debugSignals_102;
  wire [31:0] mags_0_io_debugSignals_103;
  wire [31:0] mags_0_io_debugSignals_104;
  wire [31:0] mags_0_io_debugSignals_105;
  wire [31:0] mags_0_io_debugSignals_106;
  wire [31:0] mags_0_io_debugSignals_107;
  wire [63:0] mags_0_io_TOP_AXI_AWADDR;
  wire [7:0] mags_0_io_TOP_AXI_AWLEN;
  wire  mags_0_io_TOP_AXI_AWVALID;
  wire  mags_0_io_TOP_AXI_AWREADY;
  wire  mags_0_io_TOP_AXI_ARID;
  wire [63:0] mags_0_io_TOP_AXI_ARADDR;
  wire [7:0] mags_0_io_TOP_AXI_ARLEN;
  wire [2:0] mags_0_io_TOP_AXI_ARSIZE;
  wire [1:0] mags_0_io_TOP_AXI_ARBURST;
  wire  mags_0_io_TOP_AXI_ARVALID;
  wire  mags_0_io_TOP_AXI_ARREADY;
  wire [511:0] mags_0_io_TOP_AXI_WDATA;
  wire [63:0] mags_0_io_TOP_AXI_WSTRB;
  wire  mags_0_io_TOP_AXI_WVALID;
  wire  mags_0_io_TOP_AXI_WREADY;
  wire  mags_0_io_TOP_AXI_RVALID;
  wire  mags_0_io_TOP_AXI_RREADY;
  wire  mags_0_io_TOP_AXI_BVALID;
  wire  mags_0_io_TOP_AXI_BREADY;
  wire [63:0] mags_0_io_DWIDTH_AXI_AWADDR;
  wire [7:0] mags_0_io_DWIDTH_AXI_AWLEN;
  wire  mags_0_io_DWIDTH_AXI_AWVALID;
  wire  mags_0_io_DWIDTH_AXI_AWREADY;
  wire [63:0] mags_0_io_DWIDTH_AXI_ARADDR;
  wire [7:0] mags_0_io_DWIDTH_AXI_ARLEN;
  wire [2:0] mags_0_io_DWIDTH_AXI_ARSIZE;
  wire [1:0] mags_0_io_DWIDTH_AXI_ARBURST;
  wire  mags_0_io_DWIDTH_AXI_ARVALID;
  wire  mags_0_io_DWIDTH_AXI_ARREADY;
  wire [511:0] mags_0_io_DWIDTH_AXI_WDATA;
  wire [63:0] mags_0_io_DWIDTH_AXI_WSTRB;
  wire  mags_0_io_DWIDTH_AXI_WVALID;
  wire  mags_0_io_DWIDTH_AXI_WREADY;
  wire  mags_0_io_DWIDTH_AXI_RVALID;
  wire  mags_0_io_DWIDTH_AXI_RREADY;
  wire  mags_0_io_DWIDTH_AXI_BVALID;
  wire  mags_0_io_DWIDTH_AXI_BREADY;
  wire  mags_1_clock;
  wire  mags_1_reset;
  wire  mags_1_io_enable;
  wire  mags_1_io_reset;
  wire  mags_1_io_app_loads_0_cmd_ready;
  wire  mags_1_io_app_loads_0_cmd_valid;
  wire [63:0] mags_1_io_app_loads_0_cmd_bits_addr;
  wire  mags_1_io_app_loads_0_cmd_bits_isWr;
  wire [15:0] mags_1_io_app_loads_0_cmd_bits_size;
  wire  mags_1_io_app_loads_0_rdata_ready;
  wire  mags_1_io_app_loads_0_rdata_valid;
  wire [31:0] mags_1_io_app_loads_0_rdata_bits_0;
  wire  mags_1_io_dram_cmd_ready;
  wire  mags_1_io_dram_cmd_valid;
  wire [63:0] mags_1_io_dram_cmd_bits_addr;
  wire [31:0] mags_1_io_dram_cmd_bits_size;
  wire  mags_1_io_dram_cmd_bits_isWr;
  wire [25:0] mags_1_io_dram_cmd_bits_tag_uid;
  wire [5:0] mags_1_io_dram_cmd_bits_tag_streamId;
  wire  mags_1_io_dram_wdata_ready;
  wire  mags_1_io_dram_wdata_valid;
  wire [31:0] mags_1_io_dram_wdata_bits_wdata_0;
  wire [31:0] mags_1_io_dram_wdata_bits_wdata_1;
  wire [31:0] mags_1_io_dram_wdata_bits_wdata_2;
  wire [31:0] mags_1_io_dram_wdata_bits_wdata_3;
  wire [31:0] mags_1_io_dram_wdata_bits_wdata_4;
  wire [31:0] mags_1_io_dram_wdata_bits_wdata_5;
  wire [31:0] mags_1_io_dram_wdata_bits_wdata_6;
  wire [31:0] mags_1_io_dram_wdata_bits_wdata_7;
  wire [31:0] mags_1_io_dram_wdata_bits_wdata_8;
  wire [31:0] mags_1_io_dram_wdata_bits_wdata_9;
  wire [31:0] mags_1_io_dram_wdata_bits_wdata_10;
  wire [31:0] mags_1_io_dram_wdata_bits_wdata_11;
  wire [31:0] mags_1_io_dram_wdata_bits_wdata_12;
  wire [31:0] mags_1_io_dram_wdata_bits_wdata_13;
  wire [31:0] mags_1_io_dram_wdata_bits_wdata_14;
  wire [31:0] mags_1_io_dram_wdata_bits_wdata_15;
  wire  mags_1_io_dram_wdata_bits_wstrb_0;
  wire  mags_1_io_dram_wdata_bits_wstrb_1;
  wire  mags_1_io_dram_wdata_bits_wstrb_2;
  wire  mags_1_io_dram_wdata_bits_wstrb_3;
  wire  mags_1_io_dram_wdata_bits_wstrb_4;
  wire  mags_1_io_dram_wdata_bits_wstrb_5;
  wire  mags_1_io_dram_wdata_bits_wstrb_6;
  wire  mags_1_io_dram_wdata_bits_wstrb_7;
  wire  mags_1_io_dram_wdata_bits_wstrb_8;
  wire  mags_1_io_dram_wdata_bits_wstrb_9;
  wire  mags_1_io_dram_wdata_bits_wstrb_10;
  wire  mags_1_io_dram_wdata_bits_wstrb_11;
  wire  mags_1_io_dram_wdata_bits_wstrb_12;
  wire  mags_1_io_dram_wdata_bits_wstrb_13;
  wire  mags_1_io_dram_wdata_bits_wstrb_14;
  wire  mags_1_io_dram_wdata_bits_wstrb_15;
  wire  mags_1_io_dram_wdata_bits_wstrb_16;
  wire  mags_1_io_dram_wdata_bits_wstrb_17;
  wire  mags_1_io_dram_wdata_bits_wstrb_18;
  wire  mags_1_io_dram_wdata_bits_wstrb_19;
  wire  mags_1_io_dram_wdata_bits_wstrb_20;
  wire  mags_1_io_dram_wdata_bits_wstrb_21;
  wire  mags_1_io_dram_wdata_bits_wstrb_22;
  wire  mags_1_io_dram_wdata_bits_wstrb_23;
  wire  mags_1_io_dram_wdata_bits_wstrb_24;
  wire  mags_1_io_dram_wdata_bits_wstrb_25;
  wire  mags_1_io_dram_wdata_bits_wstrb_26;
  wire  mags_1_io_dram_wdata_bits_wstrb_27;
  wire  mags_1_io_dram_wdata_bits_wstrb_28;
  wire  mags_1_io_dram_wdata_bits_wstrb_29;
  wire  mags_1_io_dram_wdata_bits_wstrb_30;
  wire  mags_1_io_dram_wdata_bits_wstrb_31;
  wire  mags_1_io_dram_wdata_bits_wstrb_32;
  wire  mags_1_io_dram_wdata_bits_wstrb_33;
  wire  mags_1_io_dram_wdata_bits_wstrb_34;
  wire  mags_1_io_dram_wdata_bits_wstrb_35;
  wire  mags_1_io_dram_wdata_bits_wstrb_36;
  wire  mags_1_io_dram_wdata_bits_wstrb_37;
  wire  mags_1_io_dram_wdata_bits_wstrb_38;
  wire  mags_1_io_dram_wdata_bits_wstrb_39;
  wire  mags_1_io_dram_wdata_bits_wstrb_40;
  wire  mags_1_io_dram_wdata_bits_wstrb_41;
  wire  mags_1_io_dram_wdata_bits_wstrb_42;
  wire  mags_1_io_dram_wdata_bits_wstrb_43;
  wire  mags_1_io_dram_wdata_bits_wstrb_44;
  wire  mags_1_io_dram_wdata_bits_wstrb_45;
  wire  mags_1_io_dram_wdata_bits_wstrb_46;
  wire  mags_1_io_dram_wdata_bits_wstrb_47;
  wire  mags_1_io_dram_wdata_bits_wstrb_48;
  wire  mags_1_io_dram_wdata_bits_wstrb_49;
  wire  mags_1_io_dram_wdata_bits_wstrb_50;
  wire  mags_1_io_dram_wdata_bits_wstrb_51;
  wire  mags_1_io_dram_wdata_bits_wstrb_52;
  wire  mags_1_io_dram_wdata_bits_wstrb_53;
  wire  mags_1_io_dram_wdata_bits_wstrb_54;
  wire  mags_1_io_dram_wdata_bits_wstrb_55;
  wire  mags_1_io_dram_wdata_bits_wstrb_56;
  wire  mags_1_io_dram_wdata_bits_wstrb_57;
  wire  mags_1_io_dram_wdata_bits_wstrb_58;
  wire  mags_1_io_dram_wdata_bits_wstrb_59;
  wire  mags_1_io_dram_wdata_bits_wstrb_60;
  wire  mags_1_io_dram_wdata_bits_wstrb_61;
  wire  mags_1_io_dram_wdata_bits_wstrb_62;
  wire  mags_1_io_dram_wdata_bits_wstrb_63;
  wire  mags_1_io_dram_rresp_ready;
  wire  mags_1_io_dram_rresp_valid;
  wire [31:0] mags_1_io_dram_rresp_bits_rdata_0;
  wire [31:0] mags_1_io_dram_rresp_bits_rdata_1;
  wire [31:0] mags_1_io_dram_rresp_bits_rdata_2;
  wire [31:0] mags_1_io_dram_rresp_bits_rdata_3;
  wire [31:0] mags_1_io_dram_rresp_bits_rdata_4;
  wire [31:0] mags_1_io_dram_rresp_bits_rdata_5;
  wire [31:0] mags_1_io_dram_rresp_bits_rdata_6;
  wire [31:0] mags_1_io_dram_rresp_bits_rdata_7;
  wire [31:0] mags_1_io_dram_rresp_bits_rdata_8;
  wire [31:0] mags_1_io_dram_rresp_bits_rdata_9;
  wire [31:0] mags_1_io_dram_rresp_bits_rdata_10;
  wire [31:0] mags_1_io_dram_rresp_bits_rdata_11;
  wire [31:0] mags_1_io_dram_rresp_bits_rdata_12;
  wire [31:0] mags_1_io_dram_rresp_bits_rdata_13;
  wire [31:0] mags_1_io_dram_rresp_bits_rdata_14;
  wire [31:0] mags_1_io_dram_rresp_bits_rdata_15;
  wire [5:0] mags_1_io_dram_rresp_bits_tag_streamId;
  wire  mags_1_io_dram_wresp_ready;
  wire  mags_1_io_dram_wresp_valid;
  wire [5:0] mags_1_io_dram_wresp_bits_tag_streamId;
  wire  mags_2_clock;
  wire  mags_2_reset;
  wire  mags_2_io_enable;
  wire  mags_2_io_reset;
  wire  mags_2_io_app_loads_0_cmd_ready;
  wire  mags_2_io_app_loads_0_cmd_valid;
  wire [63:0] mags_2_io_app_loads_0_cmd_bits_addr;
  wire  mags_2_io_app_loads_0_cmd_bits_isWr;
  wire [15:0] mags_2_io_app_loads_0_cmd_bits_size;
  wire  mags_2_io_app_loads_0_rdata_ready;
  wire  mags_2_io_app_loads_0_rdata_valid;
  wire [31:0] mags_2_io_app_loads_0_rdata_bits_0;
  wire  mags_2_io_dram_cmd_ready;
  wire  mags_2_io_dram_cmd_valid;
  wire [63:0] mags_2_io_dram_cmd_bits_addr;
  wire [31:0] mags_2_io_dram_cmd_bits_size;
  wire  mags_2_io_dram_cmd_bits_isWr;
  wire [25:0] mags_2_io_dram_cmd_bits_tag_uid;
  wire [5:0] mags_2_io_dram_cmd_bits_tag_streamId;
  wire  mags_2_io_dram_wdata_ready;
  wire  mags_2_io_dram_wdata_valid;
  wire [31:0] mags_2_io_dram_wdata_bits_wdata_0;
  wire [31:0] mags_2_io_dram_wdata_bits_wdata_1;
  wire [31:0] mags_2_io_dram_wdata_bits_wdata_2;
  wire [31:0] mags_2_io_dram_wdata_bits_wdata_3;
  wire [31:0] mags_2_io_dram_wdata_bits_wdata_4;
  wire [31:0] mags_2_io_dram_wdata_bits_wdata_5;
  wire [31:0] mags_2_io_dram_wdata_bits_wdata_6;
  wire [31:0] mags_2_io_dram_wdata_bits_wdata_7;
  wire [31:0] mags_2_io_dram_wdata_bits_wdata_8;
  wire [31:0] mags_2_io_dram_wdata_bits_wdata_9;
  wire [31:0] mags_2_io_dram_wdata_bits_wdata_10;
  wire [31:0] mags_2_io_dram_wdata_bits_wdata_11;
  wire [31:0] mags_2_io_dram_wdata_bits_wdata_12;
  wire [31:0] mags_2_io_dram_wdata_bits_wdata_13;
  wire [31:0] mags_2_io_dram_wdata_bits_wdata_14;
  wire [31:0] mags_2_io_dram_wdata_bits_wdata_15;
  wire  mags_2_io_dram_wdata_bits_wstrb_0;
  wire  mags_2_io_dram_wdata_bits_wstrb_1;
  wire  mags_2_io_dram_wdata_bits_wstrb_2;
  wire  mags_2_io_dram_wdata_bits_wstrb_3;
  wire  mags_2_io_dram_wdata_bits_wstrb_4;
  wire  mags_2_io_dram_wdata_bits_wstrb_5;
  wire  mags_2_io_dram_wdata_bits_wstrb_6;
  wire  mags_2_io_dram_wdata_bits_wstrb_7;
  wire  mags_2_io_dram_wdata_bits_wstrb_8;
  wire  mags_2_io_dram_wdata_bits_wstrb_9;
  wire  mags_2_io_dram_wdata_bits_wstrb_10;
  wire  mags_2_io_dram_wdata_bits_wstrb_11;
  wire  mags_2_io_dram_wdata_bits_wstrb_12;
  wire  mags_2_io_dram_wdata_bits_wstrb_13;
  wire  mags_2_io_dram_wdata_bits_wstrb_14;
  wire  mags_2_io_dram_wdata_bits_wstrb_15;
  wire  mags_2_io_dram_wdata_bits_wstrb_16;
  wire  mags_2_io_dram_wdata_bits_wstrb_17;
  wire  mags_2_io_dram_wdata_bits_wstrb_18;
  wire  mags_2_io_dram_wdata_bits_wstrb_19;
  wire  mags_2_io_dram_wdata_bits_wstrb_20;
  wire  mags_2_io_dram_wdata_bits_wstrb_21;
  wire  mags_2_io_dram_wdata_bits_wstrb_22;
  wire  mags_2_io_dram_wdata_bits_wstrb_23;
  wire  mags_2_io_dram_wdata_bits_wstrb_24;
  wire  mags_2_io_dram_wdata_bits_wstrb_25;
  wire  mags_2_io_dram_wdata_bits_wstrb_26;
  wire  mags_2_io_dram_wdata_bits_wstrb_27;
  wire  mags_2_io_dram_wdata_bits_wstrb_28;
  wire  mags_2_io_dram_wdata_bits_wstrb_29;
  wire  mags_2_io_dram_wdata_bits_wstrb_30;
  wire  mags_2_io_dram_wdata_bits_wstrb_31;
  wire  mags_2_io_dram_wdata_bits_wstrb_32;
  wire  mags_2_io_dram_wdata_bits_wstrb_33;
  wire  mags_2_io_dram_wdata_bits_wstrb_34;
  wire  mags_2_io_dram_wdata_bits_wstrb_35;
  wire  mags_2_io_dram_wdata_bits_wstrb_36;
  wire  mags_2_io_dram_wdata_bits_wstrb_37;
  wire  mags_2_io_dram_wdata_bits_wstrb_38;
  wire  mags_2_io_dram_wdata_bits_wstrb_39;
  wire  mags_2_io_dram_wdata_bits_wstrb_40;
  wire  mags_2_io_dram_wdata_bits_wstrb_41;
  wire  mags_2_io_dram_wdata_bits_wstrb_42;
  wire  mags_2_io_dram_wdata_bits_wstrb_43;
  wire  mags_2_io_dram_wdata_bits_wstrb_44;
  wire  mags_2_io_dram_wdata_bits_wstrb_45;
  wire  mags_2_io_dram_wdata_bits_wstrb_46;
  wire  mags_2_io_dram_wdata_bits_wstrb_47;
  wire  mags_2_io_dram_wdata_bits_wstrb_48;
  wire  mags_2_io_dram_wdata_bits_wstrb_49;
  wire  mags_2_io_dram_wdata_bits_wstrb_50;
  wire  mags_2_io_dram_wdata_bits_wstrb_51;
  wire  mags_2_io_dram_wdata_bits_wstrb_52;
  wire  mags_2_io_dram_wdata_bits_wstrb_53;
  wire  mags_2_io_dram_wdata_bits_wstrb_54;
  wire  mags_2_io_dram_wdata_bits_wstrb_55;
  wire  mags_2_io_dram_wdata_bits_wstrb_56;
  wire  mags_2_io_dram_wdata_bits_wstrb_57;
  wire  mags_2_io_dram_wdata_bits_wstrb_58;
  wire  mags_2_io_dram_wdata_bits_wstrb_59;
  wire  mags_2_io_dram_wdata_bits_wstrb_60;
  wire  mags_2_io_dram_wdata_bits_wstrb_61;
  wire  mags_2_io_dram_wdata_bits_wstrb_62;
  wire  mags_2_io_dram_wdata_bits_wstrb_63;
  wire  mags_2_io_dram_rresp_ready;
  wire  mags_2_io_dram_rresp_valid;
  wire [31:0] mags_2_io_dram_rresp_bits_rdata_0;
  wire [31:0] mags_2_io_dram_rresp_bits_rdata_1;
  wire [31:0] mags_2_io_dram_rresp_bits_rdata_2;
  wire [31:0] mags_2_io_dram_rresp_bits_rdata_3;
  wire [31:0] mags_2_io_dram_rresp_bits_rdata_4;
  wire [31:0] mags_2_io_dram_rresp_bits_rdata_5;
  wire [31:0] mags_2_io_dram_rresp_bits_rdata_6;
  wire [31:0] mags_2_io_dram_rresp_bits_rdata_7;
  wire [31:0] mags_2_io_dram_rresp_bits_rdata_8;
  wire [31:0] mags_2_io_dram_rresp_bits_rdata_9;
  wire [31:0] mags_2_io_dram_rresp_bits_rdata_10;
  wire [31:0] mags_2_io_dram_rresp_bits_rdata_11;
  wire [31:0] mags_2_io_dram_rresp_bits_rdata_12;
  wire [31:0] mags_2_io_dram_rresp_bits_rdata_13;
  wire [31:0] mags_2_io_dram_rresp_bits_rdata_14;
  wire [31:0] mags_2_io_dram_rresp_bits_rdata_15;
  wire [5:0] mags_2_io_dram_rresp_bits_tag_streamId;
  wire  mags_2_io_dram_wresp_ready;
  wire  mags_2_io_dram_wresp_valid;
  wire [5:0] mags_2_io_dram_wresp_bits_tag_streamId;
  wire  mags_3_clock;
  wire  mags_3_reset;
  wire  mags_3_io_enable;
  wire  mags_3_io_reset;
  wire  mags_3_io_app_loads_0_cmd_ready;
  wire  mags_3_io_app_loads_0_cmd_valid;
  wire [63:0] mags_3_io_app_loads_0_cmd_bits_addr;
  wire  mags_3_io_app_loads_0_cmd_bits_isWr;
  wire [15:0] mags_3_io_app_loads_0_cmd_bits_size;
  wire  mags_3_io_app_loads_0_rdata_ready;
  wire  mags_3_io_app_loads_0_rdata_valid;
  wire [31:0] mags_3_io_app_loads_0_rdata_bits_0;
  wire  mags_3_io_dram_cmd_ready;
  wire  mags_3_io_dram_cmd_valid;
  wire [63:0] mags_3_io_dram_cmd_bits_addr;
  wire [31:0] mags_3_io_dram_cmd_bits_size;
  wire  mags_3_io_dram_cmd_bits_isWr;
  wire [25:0] mags_3_io_dram_cmd_bits_tag_uid;
  wire [5:0] mags_3_io_dram_cmd_bits_tag_streamId;
  wire  mags_3_io_dram_wdata_ready;
  wire  mags_3_io_dram_wdata_valid;
  wire [31:0] mags_3_io_dram_wdata_bits_wdata_0;
  wire [31:0] mags_3_io_dram_wdata_bits_wdata_1;
  wire [31:0] mags_3_io_dram_wdata_bits_wdata_2;
  wire [31:0] mags_3_io_dram_wdata_bits_wdata_3;
  wire [31:0] mags_3_io_dram_wdata_bits_wdata_4;
  wire [31:0] mags_3_io_dram_wdata_bits_wdata_5;
  wire [31:0] mags_3_io_dram_wdata_bits_wdata_6;
  wire [31:0] mags_3_io_dram_wdata_bits_wdata_7;
  wire [31:0] mags_3_io_dram_wdata_bits_wdata_8;
  wire [31:0] mags_3_io_dram_wdata_bits_wdata_9;
  wire [31:0] mags_3_io_dram_wdata_bits_wdata_10;
  wire [31:0] mags_3_io_dram_wdata_bits_wdata_11;
  wire [31:0] mags_3_io_dram_wdata_bits_wdata_12;
  wire [31:0] mags_3_io_dram_wdata_bits_wdata_13;
  wire [31:0] mags_3_io_dram_wdata_bits_wdata_14;
  wire [31:0] mags_3_io_dram_wdata_bits_wdata_15;
  wire  mags_3_io_dram_wdata_bits_wstrb_0;
  wire  mags_3_io_dram_wdata_bits_wstrb_1;
  wire  mags_3_io_dram_wdata_bits_wstrb_2;
  wire  mags_3_io_dram_wdata_bits_wstrb_3;
  wire  mags_3_io_dram_wdata_bits_wstrb_4;
  wire  mags_3_io_dram_wdata_bits_wstrb_5;
  wire  mags_3_io_dram_wdata_bits_wstrb_6;
  wire  mags_3_io_dram_wdata_bits_wstrb_7;
  wire  mags_3_io_dram_wdata_bits_wstrb_8;
  wire  mags_3_io_dram_wdata_bits_wstrb_9;
  wire  mags_3_io_dram_wdata_bits_wstrb_10;
  wire  mags_3_io_dram_wdata_bits_wstrb_11;
  wire  mags_3_io_dram_wdata_bits_wstrb_12;
  wire  mags_3_io_dram_wdata_bits_wstrb_13;
  wire  mags_3_io_dram_wdata_bits_wstrb_14;
  wire  mags_3_io_dram_wdata_bits_wstrb_15;
  wire  mags_3_io_dram_wdata_bits_wstrb_16;
  wire  mags_3_io_dram_wdata_bits_wstrb_17;
  wire  mags_3_io_dram_wdata_bits_wstrb_18;
  wire  mags_3_io_dram_wdata_bits_wstrb_19;
  wire  mags_3_io_dram_wdata_bits_wstrb_20;
  wire  mags_3_io_dram_wdata_bits_wstrb_21;
  wire  mags_3_io_dram_wdata_bits_wstrb_22;
  wire  mags_3_io_dram_wdata_bits_wstrb_23;
  wire  mags_3_io_dram_wdata_bits_wstrb_24;
  wire  mags_3_io_dram_wdata_bits_wstrb_25;
  wire  mags_3_io_dram_wdata_bits_wstrb_26;
  wire  mags_3_io_dram_wdata_bits_wstrb_27;
  wire  mags_3_io_dram_wdata_bits_wstrb_28;
  wire  mags_3_io_dram_wdata_bits_wstrb_29;
  wire  mags_3_io_dram_wdata_bits_wstrb_30;
  wire  mags_3_io_dram_wdata_bits_wstrb_31;
  wire  mags_3_io_dram_wdata_bits_wstrb_32;
  wire  mags_3_io_dram_wdata_bits_wstrb_33;
  wire  mags_3_io_dram_wdata_bits_wstrb_34;
  wire  mags_3_io_dram_wdata_bits_wstrb_35;
  wire  mags_3_io_dram_wdata_bits_wstrb_36;
  wire  mags_3_io_dram_wdata_bits_wstrb_37;
  wire  mags_3_io_dram_wdata_bits_wstrb_38;
  wire  mags_3_io_dram_wdata_bits_wstrb_39;
  wire  mags_3_io_dram_wdata_bits_wstrb_40;
  wire  mags_3_io_dram_wdata_bits_wstrb_41;
  wire  mags_3_io_dram_wdata_bits_wstrb_42;
  wire  mags_3_io_dram_wdata_bits_wstrb_43;
  wire  mags_3_io_dram_wdata_bits_wstrb_44;
  wire  mags_3_io_dram_wdata_bits_wstrb_45;
  wire  mags_3_io_dram_wdata_bits_wstrb_46;
  wire  mags_3_io_dram_wdata_bits_wstrb_47;
  wire  mags_3_io_dram_wdata_bits_wstrb_48;
  wire  mags_3_io_dram_wdata_bits_wstrb_49;
  wire  mags_3_io_dram_wdata_bits_wstrb_50;
  wire  mags_3_io_dram_wdata_bits_wstrb_51;
  wire  mags_3_io_dram_wdata_bits_wstrb_52;
  wire  mags_3_io_dram_wdata_bits_wstrb_53;
  wire  mags_3_io_dram_wdata_bits_wstrb_54;
  wire  mags_3_io_dram_wdata_bits_wstrb_55;
  wire  mags_3_io_dram_wdata_bits_wstrb_56;
  wire  mags_3_io_dram_wdata_bits_wstrb_57;
  wire  mags_3_io_dram_wdata_bits_wstrb_58;
  wire  mags_3_io_dram_wdata_bits_wstrb_59;
  wire  mags_3_io_dram_wdata_bits_wstrb_60;
  wire  mags_3_io_dram_wdata_bits_wstrb_61;
  wire  mags_3_io_dram_wdata_bits_wstrb_62;
  wire  mags_3_io_dram_wdata_bits_wstrb_63;
  wire  mags_3_io_dram_rresp_ready;
  wire  mags_3_io_dram_rresp_valid;
  wire [31:0] mags_3_io_dram_rresp_bits_rdata_0;
  wire [31:0] mags_3_io_dram_rresp_bits_rdata_1;
  wire [31:0] mags_3_io_dram_rresp_bits_rdata_2;
  wire [31:0] mags_3_io_dram_rresp_bits_rdata_3;
  wire [31:0] mags_3_io_dram_rresp_bits_rdata_4;
  wire [31:0] mags_3_io_dram_rresp_bits_rdata_5;
  wire [31:0] mags_3_io_dram_rresp_bits_rdata_6;
  wire [31:0] mags_3_io_dram_rresp_bits_rdata_7;
  wire [31:0] mags_3_io_dram_rresp_bits_rdata_8;
  wire [31:0] mags_3_io_dram_rresp_bits_rdata_9;
  wire [31:0] mags_3_io_dram_rresp_bits_rdata_10;
  wire [31:0] mags_3_io_dram_rresp_bits_rdata_11;
  wire [31:0] mags_3_io_dram_rresp_bits_rdata_12;
  wire [31:0] mags_3_io_dram_rresp_bits_rdata_13;
  wire [31:0] mags_3_io_dram_rresp_bits_rdata_14;
  wire [31:0] mags_3_io_dram_rresp_bits_rdata_15;
  wire [5:0] mags_3_io_dram_rresp_bits_tag_streamId;
  wire  mags_3_io_dram_wresp_ready;
  wire  mags_3_io_dram_wresp_valid;
  wire [5:0] mags_3_io_dram_wresp_bits_tag_streamId;
  wire  regs_clock;
  wire  regs_reset;
  wire [31:0] regs_io_raddr;
  wire  regs_io_wen;
  wire [31:0] regs_io_waddr;
  wire [63:0] regs_io_wdata;
  wire [63:0] regs_io_rdata;
  wire  regs_io_reset;
  wire [63:0] regs_io_argIns_0;
  wire [63:0] regs_io_argIns_1;
  wire [63:0] regs_io_argIns_2;
  wire [63:0] regs_io_argIns_3;
  wire [63:0] regs_io_argIns_4;
  wire  regs_io_argOuts_0_valid;
  wire [63:0] regs_io_argOuts_0_bits;
  wire  regs_io_argOuts_1_valid;
  wire [63:0] regs_io_argOuts_1_bits;
  wire [63:0] regs_io_argOuts_2_bits;
  wire [63:0] regs_io_argOuts_3_bits;
  wire [63:0] regs_io_argOuts_4_bits;
  wire [63:0] regs_io_argOuts_5_bits;
  wire [63:0] regs_io_argOuts_6_bits;
  wire [63:0] regs_io_argOuts_7_bits;
  wire [63:0] regs_io_argOuts_8_bits;
  wire [63:0] regs_io_argOuts_9_bits;
  wire [63:0] regs_io_argOuts_10_bits;
  wire [63:0] regs_io_argOuts_11_bits;
  wire [63:0] regs_io_argOuts_12_bits;
  wire [63:0] regs_io_argOuts_13_bits;
  wire [63:0] regs_io_argOuts_14_bits;
  wire [63:0] regs_io_argOuts_15_bits;
  wire [63:0] regs_io_argOuts_16_bits;
  wire [63:0] regs_io_argOuts_17_bits;
  wire [63:0] regs_io_argOuts_18_bits;
  wire [63:0] regs_io_argOuts_19_bits;
  wire [63:0] regs_io_argOuts_20_bits;
  wire [63:0] regs_io_argOuts_21_bits;
  wire [63:0] regs_io_argOuts_22_bits;
  wire [63:0] regs_io_argOuts_23_bits;
  wire [63:0] regs_io_argOuts_24_bits;
  wire [63:0] regs_io_argOuts_25_bits;
  wire [63:0] regs_io_argOuts_26_bits;
  wire [63:0] regs_io_argOuts_27_bits;
  wire [63:0] regs_io_argOuts_28_bits;
  wire [63:0] regs_io_argOuts_29_bits;
  wire [63:0] regs_io_argOuts_30_bits;
  wire [63:0] regs_io_argOuts_31_bits;
  wire [63:0] regs_io_argOuts_32_bits;
  wire [63:0] regs_io_argOuts_33_bits;
  wire [63:0] regs_io_argOuts_34_bits;
  wire [63:0] regs_io_argOuts_35_bits;
  wire [63:0] regs_io_argOuts_36_bits;
  wire [63:0] regs_io_argOuts_37_bits;
  wire [63:0] regs_io_argOuts_38_bits;
  wire [63:0] regs_io_argOuts_39_bits;
  wire [63:0] regs_io_argOuts_40_bits;
  wire [63:0] regs_io_argOuts_41_bits;
  wire [63:0] regs_io_argOuts_42_bits;
  wire [63:0] regs_io_argOuts_43_bits;
  wire [63:0] regs_io_argOuts_44_bits;
  wire [63:0] regs_io_argOuts_45_bits;
  wire [63:0] regs_io_argOuts_46_bits;
  wire [63:0] regs_io_argOuts_47_bits;
  wire [63:0] regs_io_argOuts_48_bits;
  wire [63:0] regs_io_argOuts_49_bits;
  wire [63:0] regs_io_argOuts_50_bits;
  wire [63:0] regs_io_argOuts_51_bits;
  wire [63:0] regs_io_argOuts_52_bits;
  wire [63:0] regs_io_argOuts_53_bits;
  wire [63:0] regs_io_argOuts_54_bits;
  wire [63:0] regs_io_argOuts_55_bits;
  wire [63:0] regs_io_argOuts_56_bits;
  wire [63:0] regs_io_argOuts_57_bits;
  wire [63:0] regs_io_argOuts_58_bits;
  wire [63:0] regs_io_argOuts_59_bits;
  wire [63:0] regs_io_argOuts_60_bits;
  wire [63:0] regs_io_argOuts_61_bits;
  wire [63:0] regs_io_argOuts_62_bits;
  wire [63:0] regs_io_argOuts_63_bits;
  wire [63:0] regs_io_argOuts_64_bits;
  wire [63:0] regs_io_argOuts_65_bits;
  wire [63:0] regs_io_argOuts_66_bits;
  wire [63:0] regs_io_argOuts_67_bits;
  wire [63:0] regs_io_argOuts_68_bits;
  wire [63:0] regs_io_argOuts_69_bits;
  wire [63:0] regs_io_argOuts_70_bits;
  wire [63:0] regs_io_argOuts_71_bits;
  wire [63:0] regs_io_argOuts_72_bits;
  wire [63:0] regs_io_argOuts_73_bits;
  wire [63:0] regs_io_argOuts_74_bits;
  wire [63:0] regs_io_argOuts_75_bits;
  wire [63:0] regs_io_argOuts_76_bits;
  wire [63:0] regs_io_argOuts_77_bits;
  wire [63:0] regs_io_argOuts_78_bits;
  wire [63:0] regs_io_argOuts_79_bits;
  wire [63:0] regs_io_argOuts_80_bits;
  wire [63:0] regs_io_argOuts_81_bits;
  wire [63:0] regs_io_argOuts_82_bits;
  wire [63:0] regs_io_argOuts_83_bits;
  wire [63:0] regs_io_argOuts_84_bits;
  wire [63:0] regs_io_argOuts_85_bits;
  wire [63:0] regs_io_argOuts_86_bits;
  wire [63:0] regs_io_argOuts_87_bits;
  wire [63:0] regs_io_argOuts_88_bits;
  wire [63:0] regs_io_argOuts_89_bits;
  wire [63:0] regs_io_argOuts_90_bits;
  wire [63:0] regs_io_argOuts_91_bits;
  wire [63:0] regs_io_argOuts_92_bits;
  wire [63:0] regs_io_argOuts_93_bits;
  wire [63:0] regs_io_argOuts_94_bits;
  wire [63:0] regs_io_argOuts_95_bits;
  wire [63:0] regs_io_argOuts_96_bits;
  wire [63:0] regs_io_argOuts_97_bits;
  wire [63:0] regs_io_argOuts_98_bits;
  wire [63:0] regs_io_argOuts_99_bits;
  wire [63:0] regs_io_argOuts_100_bits;
  wire [63:0] regs_io_argOuts_101_bits;
  wire [63:0] regs_io_argOuts_102_bits;
  wire [63:0] regs_io_argOuts_103_bits;
  wire [63:0] regs_io_argOuts_104_bits;
  wire [63:0] regs_io_argOuts_105_bits;
  wire [63:0] regs_io_argOuts_106_bits;
  wire [63:0] regs_io_argOuts_107_bits;
  wire [63:0] regs_io_argOuts_108_bits;
  wire [63:0] regs_io_argOuts_109_bits;
  wire  _T_712;
  wire  _T_715;
  wire  _T_716;
  wire  localEnable;
  wire  _T_717;
  wire  localReset;
  wire  timeoutCtr_clock;
  wire  timeoutCtr_reset;
  wire  timeoutCtr_io_enable;
  wire  timeoutCtr_io_done;
  wire  depulser_clock;
  wire  depulser_reset;
  wire  depulser_io_in;
  wire  depulser_io_rst;
  wire  depulser_io_out;
  wire  _T_726;
  wire [63:0] _T_727;
  wire  status_valid;
  wire [63:0] status_bits;
  wire  _T_737;
  wire  _T_739;
  wire [1:0] _T_740;
  MAGCore mags_0 (
    .clock(mags_0_clock),
    .reset(mags_0_reset),
    .io_enable(mags_0_io_enable),
    .io_reset(mags_0_io_reset),
    .io_app_loads_0_cmd_ready(mags_0_io_app_loads_0_cmd_ready),
    .io_app_loads_0_cmd_valid(mags_0_io_app_loads_0_cmd_valid),
    .io_app_loads_0_cmd_bits_addr(mags_0_io_app_loads_0_cmd_bits_addr),
    .io_app_loads_0_cmd_bits_isWr(mags_0_io_app_loads_0_cmd_bits_isWr),
    .io_app_loads_0_cmd_bits_size(mags_0_io_app_loads_0_cmd_bits_size),
    .io_app_loads_0_rdata_ready(mags_0_io_app_loads_0_rdata_ready),
    .io_app_loads_0_rdata_valid(mags_0_io_app_loads_0_rdata_valid),
    .io_app_loads_0_rdata_bits_0(mags_0_io_app_loads_0_rdata_bits_0),
    .io_dram_cmd_ready(mags_0_io_dram_cmd_ready),
    .io_dram_cmd_valid(mags_0_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(mags_0_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(mags_0_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(mags_0_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag_uid(mags_0_io_dram_cmd_bits_tag_uid),
    .io_dram_cmd_bits_tag_streamId(mags_0_io_dram_cmd_bits_tag_streamId),
    .io_dram_wdata_ready(mags_0_io_dram_wdata_ready),
    .io_dram_wdata_valid(mags_0_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(mags_0_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(mags_0_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(mags_0_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(mags_0_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(mags_0_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(mags_0_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(mags_0_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(mags_0_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(mags_0_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(mags_0_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(mags_0_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(mags_0_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(mags_0_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(mags_0_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(mags_0_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(mags_0_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(mags_0_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(mags_0_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(mags_0_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(mags_0_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(mags_0_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(mags_0_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(mags_0_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(mags_0_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(mags_0_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(mags_0_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(mags_0_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(mags_0_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(mags_0_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(mags_0_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(mags_0_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(mags_0_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(mags_0_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(mags_0_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(mags_0_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(mags_0_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(mags_0_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(mags_0_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(mags_0_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(mags_0_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(mags_0_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(mags_0_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(mags_0_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(mags_0_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(mags_0_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(mags_0_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(mags_0_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(mags_0_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(mags_0_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(mags_0_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(mags_0_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(mags_0_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(mags_0_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(mags_0_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(mags_0_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(mags_0_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(mags_0_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(mags_0_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(mags_0_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(mags_0_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(mags_0_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(mags_0_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(mags_0_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(mags_0_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(mags_0_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(mags_0_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(mags_0_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(mags_0_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(mags_0_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(mags_0_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(mags_0_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(mags_0_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(mags_0_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(mags_0_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(mags_0_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(mags_0_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(mags_0_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(mags_0_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(mags_0_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(mags_0_io_dram_wdata_bits_wstrb_63),
    .io_dram_rresp_ready(mags_0_io_dram_rresp_ready),
    .io_dram_rresp_valid(mags_0_io_dram_rresp_valid),
    .io_dram_rresp_bits_rdata_0(mags_0_io_dram_rresp_bits_rdata_0),
    .io_dram_rresp_bits_rdata_1(mags_0_io_dram_rresp_bits_rdata_1),
    .io_dram_rresp_bits_rdata_2(mags_0_io_dram_rresp_bits_rdata_2),
    .io_dram_rresp_bits_rdata_3(mags_0_io_dram_rresp_bits_rdata_3),
    .io_dram_rresp_bits_rdata_4(mags_0_io_dram_rresp_bits_rdata_4),
    .io_dram_rresp_bits_rdata_5(mags_0_io_dram_rresp_bits_rdata_5),
    .io_dram_rresp_bits_rdata_6(mags_0_io_dram_rresp_bits_rdata_6),
    .io_dram_rresp_bits_rdata_7(mags_0_io_dram_rresp_bits_rdata_7),
    .io_dram_rresp_bits_rdata_8(mags_0_io_dram_rresp_bits_rdata_8),
    .io_dram_rresp_bits_rdata_9(mags_0_io_dram_rresp_bits_rdata_9),
    .io_dram_rresp_bits_rdata_10(mags_0_io_dram_rresp_bits_rdata_10),
    .io_dram_rresp_bits_rdata_11(mags_0_io_dram_rresp_bits_rdata_11),
    .io_dram_rresp_bits_rdata_12(mags_0_io_dram_rresp_bits_rdata_12),
    .io_dram_rresp_bits_rdata_13(mags_0_io_dram_rresp_bits_rdata_13),
    .io_dram_rresp_bits_rdata_14(mags_0_io_dram_rresp_bits_rdata_14),
    .io_dram_rresp_bits_rdata_15(mags_0_io_dram_rresp_bits_rdata_15),
    .io_dram_rresp_bits_tag_streamId(mags_0_io_dram_rresp_bits_tag_streamId),
    .io_dram_wresp_ready(mags_0_io_dram_wresp_ready),
    .io_dram_wresp_valid(mags_0_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag_streamId(mags_0_io_dram_wresp_bits_tag_streamId),
    .io_debugSignals_0(mags_0_io_debugSignals_0),
    .io_debugSignals_1(mags_0_io_debugSignals_1),
    .io_debugSignals_2(mags_0_io_debugSignals_2),
    .io_debugSignals_3(mags_0_io_debugSignals_3),
    .io_debugSignals_4(mags_0_io_debugSignals_4),
    .io_debugSignals_5(mags_0_io_debugSignals_5),
    .io_debugSignals_6(mags_0_io_debugSignals_6),
    .io_debugSignals_7(mags_0_io_debugSignals_7),
    .io_debugSignals_8(mags_0_io_debugSignals_8),
    .io_debugSignals_9(mags_0_io_debugSignals_9),
    .io_debugSignals_10(mags_0_io_debugSignals_10),
    .io_debugSignals_11(mags_0_io_debugSignals_11),
    .io_debugSignals_12(mags_0_io_debugSignals_12),
    .io_debugSignals_13(mags_0_io_debugSignals_13),
    .io_debugSignals_14(mags_0_io_debugSignals_14),
    .io_debugSignals_15(mags_0_io_debugSignals_15),
    .io_debugSignals_16(mags_0_io_debugSignals_16),
    .io_debugSignals_17(mags_0_io_debugSignals_17),
    .io_debugSignals_18(mags_0_io_debugSignals_18),
    .io_debugSignals_19(mags_0_io_debugSignals_19),
    .io_debugSignals_20(mags_0_io_debugSignals_20),
    .io_debugSignals_21(mags_0_io_debugSignals_21),
    .io_debugSignals_22(mags_0_io_debugSignals_22),
    .io_debugSignals_23(mags_0_io_debugSignals_23),
    .io_debugSignals_24(mags_0_io_debugSignals_24),
    .io_debugSignals_25(mags_0_io_debugSignals_25),
    .io_debugSignals_26(mags_0_io_debugSignals_26),
    .io_debugSignals_27(mags_0_io_debugSignals_27),
    .io_debugSignals_28(mags_0_io_debugSignals_28),
    .io_debugSignals_29(mags_0_io_debugSignals_29),
    .io_debugSignals_30(mags_0_io_debugSignals_30),
    .io_debugSignals_31(mags_0_io_debugSignals_31),
    .io_debugSignals_32(mags_0_io_debugSignals_32),
    .io_debugSignals_33(mags_0_io_debugSignals_33),
    .io_debugSignals_34(mags_0_io_debugSignals_34),
    .io_debugSignals_35(mags_0_io_debugSignals_35),
    .io_debugSignals_36(mags_0_io_debugSignals_36),
    .io_debugSignals_37(mags_0_io_debugSignals_37),
    .io_debugSignals_38(mags_0_io_debugSignals_38),
    .io_debugSignals_39(mags_0_io_debugSignals_39),
    .io_debugSignals_40(mags_0_io_debugSignals_40),
    .io_debugSignals_41(mags_0_io_debugSignals_41),
    .io_debugSignals_42(mags_0_io_debugSignals_42),
    .io_debugSignals_43(mags_0_io_debugSignals_43),
    .io_debugSignals_44(mags_0_io_debugSignals_44),
    .io_debugSignals_45(mags_0_io_debugSignals_45),
    .io_debugSignals_46(mags_0_io_debugSignals_46),
    .io_debugSignals_47(mags_0_io_debugSignals_47),
    .io_debugSignals_48(mags_0_io_debugSignals_48),
    .io_debugSignals_49(mags_0_io_debugSignals_49),
    .io_debugSignals_50(mags_0_io_debugSignals_50),
    .io_debugSignals_51(mags_0_io_debugSignals_51),
    .io_debugSignals_52(mags_0_io_debugSignals_52),
    .io_debugSignals_53(mags_0_io_debugSignals_53),
    .io_debugSignals_54(mags_0_io_debugSignals_54),
    .io_debugSignals_55(mags_0_io_debugSignals_55),
    .io_debugSignals_56(mags_0_io_debugSignals_56),
    .io_debugSignals_57(mags_0_io_debugSignals_57),
    .io_debugSignals_58(mags_0_io_debugSignals_58),
    .io_debugSignals_59(mags_0_io_debugSignals_59),
    .io_debugSignals_60(mags_0_io_debugSignals_60),
    .io_debugSignals_61(mags_0_io_debugSignals_61),
    .io_debugSignals_62(mags_0_io_debugSignals_62),
    .io_debugSignals_63(mags_0_io_debugSignals_63),
    .io_debugSignals_64(mags_0_io_debugSignals_64),
    .io_debugSignals_65(mags_0_io_debugSignals_65),
    .io_debugSignals_66(mags_0_io_debugSignals_66),
    .io_debugSignals_67(mags_0_io_debugSignals_67),
    .io_debugSignals_68(mags_0_io_debugSignals_68),
    .io_debugSignals_69(mags_0_io_debugSignals_69),
    .io_debugSignals_70(mags_0_io_debugSignals_70),
    .io_debugSignals_71(mags_0_io_debugSignals_71),
    .io_debugSignals_72(mags_0_io_debugSignals_72),
    .io_debugSignals_73(mags_0_io_debugSignals_73),
    .io_debugSignals_74(mags_0_io_debugSignals_74),
    .io_debugSignals_75(mags_0_io_debugSignals_75),
    .io_debugSignals_76(mags_0_io_debugSignals_76),
    .io_debugSignals_77(mags_0_io_debugSignals_77),
    .io_debugSignals_78(mags_0_io_debugSignals_78),
    .io_debugSignals_79(mags_0_io_debugSignals_79),
    .io_debugSignals_80(mags_0_io_debugSignals_80),
    .io_debugSignals_81(mags_0_io_debugSignals_81),
    .io_debugSignals_82(mags_0_io_debugSignals_82),
    .io_debugSignals_83(mags_0_io_debugSignals_83),
    .io_debugSignals_84(mags_0_io_debugSignals_84),
    .io_debugSignals_85(mags_0_io_debugSignals_85),
    .io_debugSignals_86(mags_0_io_debugSignals_86),
    .io_debugSignals_87(mags_0_io_debugSignals_87),
    .io_debugSignals_88(mags_0_io_debugSignals_88),
    .io_debugSignals_89(mags_0_io_debugSignals_89),
    .io_debugSignals_90(mags_0_io_debugSignals_90),
    .io_debugSignals_91(mags_0_io_debugSignals_91),
    .io_debugSignals_92(mags_0_io_debugSignals_92),
    .io_debugSignals_93(mags_0_io_debugSignals_93),
    .io_debugSignals_94(mags_0_io_debugSignals_94),
    .io_debugSignals_95(mags_0_io_debugSignals_95),
    .io_debugSignals_96(mags_0_io_debugSignals_96),
    .io_debugSignals_97(mags_0_io_debugSignals_97),
    .io_debugSignals_98(mags_0_io_debugSignals_98),
    .io_debugSignals_99(mags_0_io_debugSignals_99),
    .io_debugSignals_100(mags_0_io_debugSignals_100),
    .io_debugSignals_101(mags_0_io_debugSignals_101),
    .io_debugSignals_102(mags_0_io_debugSignals_102),
    .io_debugSignals_103(mags_0_io_debugSignals_103),
    .io_debugSignals_104(mags_0_io_debugSignals_104),
    .io_debugSignals_105(mags_0_io_debugSignals_105),
    .io_debugSignals_106(mags_0_io_debugSignals_106),
    .io_debugSignals_107(mags_0_io_debugSignals_107),
    .io_TOP_AXI_AWADDR(mags_0_io_TOP_AXI_AWADDR),
    .io_TOP_AXI_AWLEN(mags_0_io_TOP_AXI_AWLEN),
    .io_TOP_AXI_AWVALID(mags_0_io_TOP_AXI_AWVALID),
    .io_TOP_AXI_AWREADY(mags_0_io_TOP_AXI_AWREADY),
    .io_TOP_AXI_ARID(mags_0_io_TOP_AXI_ARID),
    .io_TOP_AXI_ARADDR(mags_0_io_TOP_AXI_ARADDR),
    .io_TOP_AXI_ARLEN(mags_0_io_TOP_AXI_ARLEN),
    .io_TOP_AXI_ARSIZE(mags_0_io_TOP_AXI_ARSIZE),
    .io_TOP_AXI_ARBURST(mags_0_io_TOP_AXI_ARBURST),
    .io_TOP_AXI_ARVALID(mags_0_io_TOP_AXI_ARVALID),
    .io_TOP_AXI_ARREADY(mags_0_io_TOP_AXI_ARREADY),
    .io_TOP_AXI_WDATA(mags_0_io_TOP_AXI_WDATA),
    .io_TOP_AXI_WSTRB(mags_0_io_TOP_AXI_WSTRB),
    .io_TOP_AXI_WVALID(mags_0_io_TOP_AXI_WVALID),
    .io_TOP_AXI_WREADY(mags_0_io_TOP_AXI_WREADY),
    .io_TOP_AXI_RVALID(mags_0_io_TOP_AXI_RVALID),
    .io_TOP_AXI_RREADY(mags_0_io_TOP_AXI_RREADY),
    .io_TOP_AXI_BVALID(mags_0_io_TOP_AXI_BVALID),
    .io_TOP_AXI_BREADY(mags_0_io_TOP_AXI_BREADY),
    .io_DWIDTH_AXI_AWADDR(mags_0_io_DWIDTH_AXI_AWADDR),
    .io_DWIDTH_AXI_AWLEN(mags_0_io_DWIDTH_AXI_AWLEN),
    .io_DWIDTH_AXI_AWVALID(mags_0_io_DWIDTH_AXI_AWVALID),
    .io_DWIDTH_AXI_AWREADY(mags_0_io_DWIDTH_AXI_AWREADY),
    .io_DWIDTH_AXI_ARADDR(mags_0_io_DWIDTH_AXI_ARADDR),
    .io_DWIDTH_AXI_ARLEN(mags_0_io_DWIDTH_AXI_ARLEN),
    .io_DWIDTH_AXI_ARSIZE(mags_0_io_DWIDTH_AXI_ARSIZE),
    .io_DWIDTH_AXI_ARBURST(mags_0_io_DWIDTH_AXI_ARBURST),
    .io_DWIDTH_AXI_ARVALID(mags_0_io_DWIDTH_AXI_ARVALID),
    .io_DWIDTH_AXI_ARREADY(mags_0_io_DWIDTH_AXI_ARREADY),
    .io_DWIDTH_AXI_WDATA(mags_0_io_DWIDTH_AXI_WDATA),
    .io_DWIDTH_AXI_WSTRB(mags_0_io_DWIDTH_AXI_WSTRB),
    .io_DWIDTH_AXI_WVALID(mags_0_io_DWIDTH_AXI_WVALID),
    .io_DWIDTH_AXI_WREADY(mags_0_io_DWIDTH_AXI_WREADY),
    .io_DWIDTH_AXI_RVALID(mags_0_io_DWIDTH_AXI_RVALID),
    .io_DWIDTH_AXI_RREADY(mags_0_io_DWIDTH_AXI_RREADY),
    .io_DWIDTH_AXI_BVALID(mags_0_io_DWIDTH_AXI_BVALID),
    .io_DWIDTH_AXI_BREADY(mags_0_io_DWIDTH_AXI_BREADY)
  );
  MAGCore_1 mags_1 (
    .clock(mags_1_clock),
    .reset(mags_1_reset),
    .io_enable(mags_1_io_enable),
    .io_reset(mags_1_io_reset),
    .io_app_loads_0_cmd_ready(mags_1_io_app_loads_0_cmd_ready),
    .io_app_loads_0_cmd_valid(mags_1_io_app_loads_0_cmd_valid),
    .io_app_loads_0_cmd_bits_addr(mags_1_io_app_loads_0_cmd_bits_addr),
    .io_app_loads_0_cmd_bits_isWr(mags_1_io_app_loads_0_cmd_bits_isWr),
    .io_app_loads_0_cmd_bits_size(mags_1_io_app_loads_0_cmd_bits_size),
    .io_app_loads_0_rdata_ready(mags_1_io_app_loads_0_rdata_ready),
    .io_app_loads_0_rdata_valid(mags_1_io_app_loads_0_rdata_valid),
    .io_app_loads_0_rdata_bits_0(mags_1_io_app_loads_0_rdata_bits_0),
    .io_dram_cmd_ready(mags_1_io_dram_cmd_ready),
    .io_dram_cmd_valid(mags_1_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(mags_1_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(mags_1_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(mags_1_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag_uid(mags_1_io_dram_cmd_bits_tag_uid),
    .io_dram_cmd_bits_tag_streamId(mags_1_io_dram_cmd_bits_tag_streamId),
    .io_dram_wdata_ready(mags_1_io_dram_wdata_ready),
    .io_dram_wdata_valid(mags_1_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(mags_1_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(mags_1_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(mags_1_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(mags_1_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(mags_1_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(mags_1_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(mags_1_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(mags_1_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(mags_1_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(mags_1_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(mags_1_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(mags_1_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(mags_1_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(mags_1_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(mags_1_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(mags_1_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(mags_1_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(mags_1_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(mags_1_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(mags_1_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(mags_1_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(mags_1_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(mags_1_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(mags_1_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(mags_1_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(mags_1_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(mags_1_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(mags_1_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(mags_1_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(mags_1_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(mags_1_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(mags_1_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(mags_1_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(mags_1_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(mags_1_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(mags_1_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(mags_1_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(mags_1_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(mags_1_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(mags_1_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(mags_1_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(mags_1_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(mags_1_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(mags_1_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(mags_1_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(mags_1_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(mags_1_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(mags_1_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(mags_1_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(mags_1_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(mags_1_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(mags_1_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(mags_1_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(mags_1_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(mags_1_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(mags_1_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(mags_1_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(mags_1_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(mags_1_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(mags_1_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(mags_1_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(mags_1_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(mags_1_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(mags_1_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(mags_1_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(mags_1_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(mags_1_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(mags_1_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(mags_1_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(mags_1_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(mags_1_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(mags_1_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(mags_1_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(mags_1_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(mags_1_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(mags_1_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(mags_1_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(mags_1_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(mags_1_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(mags_1_io_dram_wdata_bits_wstrb_63),
    .io_dram_rresp_ready(mags_1_io_dram_rresp_ready),
    .io_dram_rresp_valid(mags_1_io_dram_rresp_valid),
    .io_dram_rresp_bits_rdata_0(mags_1_io_dram_rresp_bits_rdata_0),
    .io_dram_rresp_bits_rdata_1(mags_1_io_dram_rresp_bits_rdata_1),
    .io_dram_rresp_bits_rdata_2(mags_1_io_dram_rresp_bits_rdata_2),
    .io_dram_rresp_bits_rdata_3(mags_1_io_dram_rresp_bits_rdata_3),
    .io_dram_rresp_bits_rdata_4(mags_1_io_dram_rresp_bits_rdata_4),
    .io_dram_rresp_bits_rdata_5(mags_1_io_dram_rresp_bits_rdata_5),
    .io_dram_rresp_bits_rdata_6(mags_1_io_dram_rresp_bits_rdata_6),
    .io_dram_rresp_bits_rdata_7(mags_1_io_dram_rresp_bits_rdata_7),
    .io_dram_rresp_bits_rdata_8(mags_1_io_dram_rresp_bits_rdata_8),
    .io_dram_rresp_bits_rdata_9(mags_1_io_dram_rresp_bits_rdata_9),
    .io_dram_rresp_bits_rdata_10(mags_1_io_dram_rresp_bits_rdata_10),
    .io_dram_rresp_bits_rdata_11(mags_1_io_dram_rresp_bits_rdata_11),
    .io_dram_rresp_bits_rdata_12(mags_1_io_dram_rresp_bits_rdata_12),
    .io_dram_rresp_bits_rdata_13(mags_1_io_dram_rresp_bits_rdata_13),
    .io_dram_rresp_bits_rdata_14(mags_1_io_dram_rresp_bits_rdata_14),
    .io_dram_rresp_bits_rdata_15(mags_1_io_dram_rresp_bits_rdata_15),
    .io_dram_rresp_bits_tag_streamId(mags_1_io_dram_rresp_bits_tag_streamId),
    .io_dram_wresp_ready(mags_1_io_dram_wresp_ready),
    .io_dram_wresp_valid(mags_1_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag_streamId(mags_1_io_dram_wresp_bits_tag_streamId)
  );
  MAGCore_1 mags_2 (
    .clock(mags_2_clock),
    .reset(mags_2_reset),
    .io_enable(mags_2_io_enable),
    .io_reset(mags_2_io_reset),
    .io_app_loads_0_cmd_ready(mags_2_io_app_loads_0_cmd_ready),
    .io_app_loads_0_cmd_valid(mags_2_io_app_loads_0_cmd_valid),
    .io_app_loads_0_cmd_bits_addr(mags_2_io_app_loads_0_cmd_bits_addr),
    .io_app_loads_0_cmd_bits_isWr(mags_2_io_app_loads_0_cmd_bits_isWr),
    .io_app_loads_0_cmd_bits_size(mags_2_io_app_loads_0_cmd_bits_size),
    .io_app_loads_0_rdata_ready(mags_2_io_app_loads_0_rdata_ready),
    .io_app_loads_0_rdata_valid(mags_2_io_app_loads_0_rdata_valid),
    .io_app_loads_0_rdata_bits_0(mags_2_io_app_loads_0_rdata_bits_0),
    .io_dram_cmd_ready(mags_2_io_dram_cmd_ready),
    .io_dram_cmd_valid(mags_2_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(mags_2_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(mags_2_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(mags_2_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag_uid(mags_2_io_dram_cmd_bits_tag_uid),
    .io_dram_cmd_bits_tag_streamId(mags_2_io_dram_cmd_bits_tag_streamId),
    .io_dram_wdata_ready(mags_2_io_dram_wdata_ready),
    .io_dram_wdata_valid(mags_2_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(mags_2_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(mags_2_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(mags_2_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(mags_2_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(mags_2_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(mags_2_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(mags_2_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(mags_2_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(mags_2_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(mags_2_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(mags_2_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(mags_2_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(mags_2_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(mags_2_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(mags_2_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(mags_2_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(mags_2_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(mags_2_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(mags_2_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(mags_2_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(mags_2_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(mags_2_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(mags_2_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(mags_2_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(mags_2_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(mags_2_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(mags_2_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(mags_2_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(mags_2_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(mags_2_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(mags_2_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(mags_2_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(mags_2_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(mags_2_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(mags_2_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(mags_2_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(mags_2_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(mags_2_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(mags_2_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(mags_2_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(mags_2_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(mags_2_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(mags_2_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(mags_2_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(mags_2_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(mags_2_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(mags_2_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(mags_2_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(mags_2_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(mags_2_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(mags_2_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(mags_2_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(mags_2_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(mags_2_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(mags_2_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(mags_2_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(mags_2_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(mags_2_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(mags_2_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(mags_2_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(mags_2_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(mags_2_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(mags_2_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(mags_2_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(mags_2_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(mags_2_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(mags_2_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(mags_2_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(mags_2_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(mags_2_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(mags_2_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(mags_2_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(mags_2_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(mags_2_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(mags_2_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(mags_2_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(mags_2_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(mags_2_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(mags_2_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(mags_2_io_dram_wdata_bits_wstrb_63),
    .io_dram_rresp_ready(mags_2_io_dram_rresp_ready),
    .io_dram_rresp_valid(mags_2_io_dram_rresp_valid),
    .io_dram_rresp_bits_rdata_0(mags_2_io_dram_rresp_bits_rdata_0),
    .io_dram_rresp_bits_rdata_1(mags_2_io_dram_rresp_bits_rdata_1),
    .io_dram_rresp_bits_rdata_2(mags_2_io_dram_rresp_bits_rdata_2),
    .io_dram_rresp_bits_rdata_3(mags_2_io_dram_rresp_bits_rdata_3),
    .io_dram_rresp_bits_rdata_4(mags_2_io_dram_rresp_bits_rdata_4),
    .io_dram_rresp_bits_rdata_5(mags_2_io_dram_rresp_bits_rdata_5),
    .io_dram_rresp_bits_rdata_6(mags_2_io_dram_rresp_bits_rdata_6),
    .io_dram_rresp_bits_rdata_7(mags_2_io_dram_rresp_bits_rdata_7),
    .io_dram_rresp_bits_rdata_8(mags_2_io_dram_rresp_bits_rdata_8),
    .io_dram_rresp_bits_rdata_9(mags_2_io_dram_rresp_bits_rdata_9),
    .io_dram_rresp_bits_rdata_10(mags_2_io_dram_rresp_bits_rdata_10),
    .io_dram_rresp_bits_rdata_11(mags_2_io_dram_rresp_bits_rdata_11),
    .io_dram_rresp_bits_rdata_12(mags_2_io_dram_rresp_bits_rdata_12),
    .io_dram_rresp_bits_rdata_13(mags_2_io_dram_rresp_bits_rdata_13),
    .io_dram_rresp_bits_rdata_14(mags_2_io_dram_rresp_bits_rdata_14),
    .io_dram_rresp_bits_rdata_15(mags_2_io_dram_rresp_bits_rdata_15),
    .io_dram_rresp_bits_tag_streamId(mags_2_io_dram_rresp_bits_tag_streamId),
    .io_dram_wresp_ready(mags_2_io_dram_wresp_ready),
    .io_dram_wresp_valid(mags_2_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag_streamId(mags_2_io_dram_wresp_bits_tag_streamId)
  );
  MAGCore_1 mags_3 (
    .clock(mags_3_clock),
    .reset(mags_3_reset),
    .io_enable(mags_3_io_enable),
    .io_reset(mags_3_io_reset),
    .io_app_loads_0_cmd_ready(mags_3_io_app_loads_0_cmd_ready),
    .io_app_loads_0_cmd_valid(mags_3_io_app_loads_0_cmd_valid),
    .io_app_loads_0_cmd_bits_addr(mags_3_io_app_loads_0_cmd_bits_addr),
    .io_app_loads_0_cmd_bits_isWr(mags_3_io_app_loads_0_cmd_bits_isWr),
    .io_app_loads_0_cmd_bits_size(mags_3_io_app_loads_0_cmd_bits_size),
    .io_app_loads_0_rdata_ready(mags_3_io_app_loads_0_rdata_ready),
    .io_app_loads_0_rdata_valid(mags_3_io_app_loads_0_rdata_valid),
    .io_app_loads_0_rdata_bits_0(mags_3_io_app_loads_0_rdata_bits_0),
    .io_dram_cmd_ready(mags_3_io_dram_cmd_ready),
    .io_dram_cmd_valid(mags_3_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(mags_3_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(mags_3_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(mags_3_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag_uid(mags_3_io_dram_cmd_bits_tag_uid),
    .io_dram_cmd_bits_tag_streamId(mags_3_io_dram_cmd_bits_tag_streamId),
    .io_dram_wdata_ready(mags_3_io_dram_wdata_ready),
    .io_dram_wdata_valid(mags_3_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(mags_3_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(mags_3_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(mags_3_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(mags_3_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(mags_3_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(mags_3_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(mags_3_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(mags_3_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(mags_3_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(mags_3_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(mags_3_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(mags_3_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(mags_3_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(mags_3_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(mags_3_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(mags_3_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(mags_3_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(mags_3_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(mags_3_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(mags_3_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(mags_3_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(mags_3_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(mags_3_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(mags_3_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(mags_3_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(mags_3_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(mags_3_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(mags_3_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(mags_3_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(mags_3_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(mags_3_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(mags_3_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(mags_3_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(mags_3_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(mags_3_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(mags_3_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(mags_3_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(mags_3_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(mags_3_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(mags_3_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(mags_3_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(mags_3_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(mags_3_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(mags_3_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(mags_3_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(mags_3_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(mags_3_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(mags_3_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(mags_3_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(mags_3_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(mags_3_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(mags_3_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(mags_3_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(mags_3_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(mags_3_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(mags_3_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(mags_3_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(mags_3_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(mags_3_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(mags_3_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(mags_3_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(mags_3_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(mags_3_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(mags_3_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(mags_3_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(mags_3_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(mags_3_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(mags_3_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(mags_3_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(mags_3_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(mags_3_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(mags_3_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(mags_3_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(mags_3_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(mags_3_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(mags_3_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(mags_3_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(mags_3_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(mags_3_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(mags_3_io_dram_wdata_bits_wstrb_63),
    .io_dram_rresp_ready(mags_3_io_dram_rresp_ready),
    .io_dram_rresp_valid(mags_3_io_dram_rresp_valid),
    .io_dram_rresp_bits_rdata_0(mags_3_io_dram_rresp_bits_rdata_0),
    .io_dram_rresp_bits_rdata_1(mags_3_io_dram_rresp_bits_rdata_1),
    .io_dram_rresp_bits_rdata_2(mags_3_io_dram_rresp_bits_rdata_2),
    .io_dram_rresp_bits_rdata_3(mags_3_io_dram_rresp_bits_rdata_3),
    .io_dram_rresp_bits_rdata_4(mags_3_io_dram_rresp_bits_rdata_4),
    .io_dram_rresp_bits_rdata_5(mags_3_io_dram_rresp_bits_rdata_5),
    .io_dram_rresp_bits_rdata_6(mags_3_io_dram_rresp_bits_rdata_6),
    .io_dram_rresp_bits_rdata_7(mags_3_io_dram_rresp_bits_rdata_7),
    .io_dram_rresp_bits_rdata_8(mags_3_io_dram_rresp_bits_rdata_8),
    .io_dram_rresp_bits_rdata_9(mags_3_io_dram_rresp_bits_rdata_9),
    .io_dram_rresp_bits_rdata_10(mags_3_io_dram_rresp_bits_rdata_10),
    .io_dram_rresp_bits_rdata_11(mags_3_io_dram_rresp_bits_rdata_11),
    .io_dram_rresp_bits_rdata_12(mags_3_io_dram_rresp_bits_rdata_12),
    .io_dram_rresp_bits_rdata_13(mags_3_io_dram_rresp_bits_rdata_13),
    .io_dram_rresp_bits_rdata_14(mags_3_io_dram_rresp_bits_rdata_14),
    .io_dram_rresp_bits_rdata_15(mags_3_io_dram_rresp_bits_rdata_15),
    .io_dram_rresp_bits_tag_streamId(mags_3_io_dram_rresp_bits_tag_streamId),
    .io_dram_wresp_ready(mags_3_io_dram_wresp_ready),
    .io_dram_wresp_valid(mags_3_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag_streamId(mags_3_io_dram_wresp_bits_tag_streamId)
  );
  RegFile regs (
    .clock(regs_clock),
    .reset(regs_reset),
    .io_raddr(regs_io_raddr),
    .io_wen(regs_io_wen),
    .io_waddr(regs_io_waddr),
    .io_wdata(regs_io_wdata),
    .io_rdata(regs_io_rdata),
    .io_reset(regs_io_reset),
    .io_argIns_0(regs_io_argIns_0),
    .io_argIns_1(regs_io_argIns_1),
    .io_argIns_2(regs_io_argIns_2),
    .io_argIns_3(regs_io_argIns_3),
    .io_argIns_4(regs_io_argIns_4),
    .io_argOuts_0_valid(regs_io_argOuts_0_valid),
    .io_argOuts_0_bits(regs_io_argOuts_0_bits),
    .io_argOuts_1_valid(regs_io_argOuts_1_valid),
    .io_argOuts_1_bits(regs_io_argOuts_1_bits),
    .io_argOuts_2_bits(regs_io_argOuts_2_bits),
    .io_argOuts_3_bits(regs_io_argOuts_3_bits),
    .io_argOuts_4_bits(regs_io_argOuts_4_bits),
    .io_argOuts_5_bits(regs_io_argOuts_5_bits),
    .io_argOuts_6_bits(regs_io_argOuts_6_bits),
    .io_argOuts_7_bits(regs_io_argOuts_7_bits),
    .io_argOuts_8_bits(regs_io_argOuts_8_bits),
    .io_argOuts_9_bits(regs_io_argOuts_9_bits),
    .io_argOuts_10_bits(regs_io_argOuts_10_bits),
    .io_argOuts_11_bits(regs_io_argOuts_11_bits),
    .io_argOuts_12_bits(regs_io_argOuts_12_bits),
    .io_argOuts_13_bits(regs_io_argOuts_13_bits),
    .io_argOuts_14_bits(regs_io_argOuts_14_bits),
    .io_argOuts_15_bits(regs_io_argOuts_15_bits),
    .io_argOuts_16_bits(regs_io_argOuts_16_bits),
    .io_argOuts_17_bits(regs_io_argOuts_17_bits),
    .io_argOuts_18_bits(regs_io_argOuts_18_bits),
    .io_argOuts_19_bits(regs_io_argOuts_19_bits),
    .io_argOuts_20_bits(regs_io_argOuts_20_bits),
    .io_argOuts_21_bits(regs_io_argOuts_21_bits),
    .io_argOuts_22_bits(regs_io_argOuts_22_bits),
    .io_argOuts_23_bits(regs_io_argOuts_23_bits),
    .io_argOuts_24_bits(regs_io_argOuts_24_bits),
    .io_argOuts_25_bits(regs_io_argOuts_25_bits),
    .io_argOuts_26_bits(regs_io_argOuts_26_bits),
    .io_argOuts_27_bits(regs_io_argOuts_27_bits),
    .io_argOuts_28_bits(regs_io_argOuts_28_bits),
    .io_argOuts_29_bits(regs_io_argOuts_29_bits),
    .io_argOuts_30_bits(regs_io_argOuts_30_bits),
    .io_argOuts_31_bits(regs_io_argOuts_31_bits),
    .io_argOuts_32_bits(regs_io_argOuts_32_bits),
    .io_argOuts_33_bits(regs_io_argOuts_33_bits),
    .io_argOuts_34_bits(regs_io_argOuts_34_bits),
    .io_argOuts_35_bits(regs_io_argOuts_35_bits),
    .io_argOuts_36_bits(regs_io_argOuts_36_bits),
    .io_argOuts_37_bits(regs_io_argOuts_37_bits),
    .io_argOuts_38_bits(regs_io_argOuts_38_bits),
    .io_argOuts_39_bits(regs_io_argOuts_39_bits),
    .io_argOuts_40_bits(regs_io_argOuts_40_bits),
    .io_argOuts_41_bits(regs_io_argOuts_41_bits),
    .io_argOuts_42_bits(regs_io_argOuts_42_bits),
    .io_argOuts_43_bits(regs_io_argOuts_43_bits),
    .io_argOuts_44_bits(regs_io_argOuts_44_bits),
    .io_argOuts_45_bits(regs_io_argOuts_45_bits),
    .io_argOuts_46_bits(regs_io_argOuts_46_bits),
    .io_argOuts_47_bits(regs_io_argOuts_47_bits),
    .io_argOuts_48_bits(regs_io_argOuts_48_bits),
    .io_argOuts_49_bits(regs_io_argOuts_49_bits),
    .io_argOuts_50_bits(regs_io_argOuts_50_bits),
    .io_argOuts_51_bits(regs_io_argOuts_51_bits),
    .io_argOuts_52_bits(regs_io_argOuts_52_bits),
    .io_argOuts_53_bits(regs_io_argOuts_53_bits),
    .io_argOuts_54_bits(regs_io_argOuts_54_bits),
    .io_argOuts_55_bits(regs_io_argOuts_55_bits),
    .io_argOuts_56_bits(regs_io_argOuts_56_bits),
    .io_argOuts_57_bits(regs_io_argOuts_57_bits),
    .io_argOuts_58_bits(regs_io_argOuts_58_bits),
    .io_argOuts_59_bits(regs_io_argOuts_59_bits),
    .io_argOuts_60_bits(regs_io_argOuts_60_bits),
    .io_argOuts_61_bits(regs_io_argOuts_61_bits),
    .io_argOuts_62_bits(regs_io_argOuts_62_bits),
    .io_argOuts_63_bits(regs_io_argOuts_63_bits),
    .io_argOuts_64_bits(regs_io_argOuts_64_bits),
    .io_argOuts_65_bits(regs_io_argOuts_65_bits),
    .io_argOuts_66_bits(regs_io_argOuts_66_bits),
    .io_argOuts_67_bits(regs_io_argOuts_67_bits),
    .io_argOuts_68_bits(regs_io_argOuts_68_bits),
    .io_argOuts_69_bits(regs_io_argOuts_69_bits),
    .io_argOuts_70_bits(regs_io_argOuts_70_bits),
    .io_argOuts_71_bits(regs_io_argOuts_71_bits),
    .io_argOuts_72_bits(regs_io_argOuts_72_bits),
    .io_argOuts_73_bits(regs_io_argOuts_73_bits),
    .io_argOuts_74_bits(regs_io_argOuts_74_bits),
    .io_argOuts_75_bits(regs_io_argOuts_75_bits),
    .io_argOuts_76_bits(regs_io_argOuts_76_bits),
    .io_argOuts_77_bits(regs_io_argOuts_77_bits),
    .io_argOuts_78_bits(regs_io_argOuts_78_bits),
    .io_argOuts_79_bits(regs_io_argOuts_79_bits),
    .io_argOuts_80_bits(regs_io_argOuts_80_bits),
    .io_argOuts_81_bits(regs_io_argOuts_81_bits),
    .io_argOuts_82_bits(regs_io_argOuts_82_bits),
    .io_argOuts_83_bits(regs_io_argOuts_83_bits),
    .io_argOuts_84_bits(regs_io_argOuts_84_bits),
    .io_argOuts_85_bits(regs_io_argOuts_85_bits),
    .io_argOuts_86_bits(regs_io_argOuts_86_bits),
    .io_argOuts_87_bits(regs_io_argOuts_87_bits),
    .io_argOuts_88_bits(regs_io_argOuts_88_bits),
    .io_argOuts_89_bits(regs_io_argOuts_89_bits),
    .io_argOuts_90_bits(regs_io_argOuts_90_bits),
    .io_argOuts_91_bits(regs_io_argOuts_91_bits),
    .io_argOuts_92_bits(regs_io_argOuts_92_bits),
    .io_argOuts_93_bits(regs_io_argOuts_93_bits),
    .io_argOuts_94_bits(regs_io_argOuts_94_bits),
    .io_argOuts_95_bits(regs_io_argOuts_95_bits),
    .io_argOuts_96_bits(regs_io_argOuts_96_bits),
    .io_argOuts_97_bits(regs_io_argOuts_97_bits),
    .io_argOuts_98_bits(regs_io_argOuts_98_bits),
    .io_argOuts_99_bits(regs_io_argOuts_99_bits),
    .io_argOuts_100_bits(regs_io_argOuts_100_bits),
    .io_argOuts_101_bits(regs_io_argOuts_101_bits),
    .io_argOuts_102_bits(regs_io_argOuts_102_bits),
    .io_argOuts_103_bits(regs_io_argOuts_103_bits),
    .io_argOuts_104_bits(regs_io_argOuts_104_bits),
    .io_argOuts_105_bits(regs_io_argOuts_105_bits),
    .io_argOuts_106_bits(regs_io_argOuts_106_bits),
    .io_argOuts_107_bits(regs_io_argOuts_107_bits),
    .io_argOuts_108_bits(regs_io_argOuts_108_bits),
    .io_argOuts_109_bits(regs_io_argOuts_109_bits)
  );
  Counter_443 timeoutCtr (
    .clock(timeoutCtr_clock),
    .reset(timeoutCtr_reset),
    .io_enable(timeoutCtr_io_enable),
    .io_done(timeoutCtr_io_done)
  );
  Depulser depulser (
    .clock(depulser_clock),
    .reset(depulser_reset),
    .io_in(depulser_io_in),
    .io_rst(depulser_io_rst),
    .io_out(depulser_io_out)
  );
  assign _T_712 = regs_io_argIns_0[0];
  assign _T_715 = regs_io_argIns_1[0];
  assign _T_716 = ~ _T_715;
  assign localEnable = _T_712 & _T_716;
  assign _T_717 = regs_io_argIns_0[1];
  assign localReset = _T_717 | reset;
  assign _T_726 = io_done | timeoutCtr_io_done;
  assign _T_727 = ~ regs_io_argIns_0;
  assign _T_737 = _T_712 & timeoutCtr_io_done;
  assign _T_739 = _T_712 & depulser_io_out;
  assign _T_740 = {_T_737,_T_739};
  assign io_rdata = regs_io_rdata;
  assign io_enable = localEnable;
  assign io_reset = localReset;
  assign io_argIns_0 = regs_io_argIns_2;
  assign io_argIns_1 = regs_io_argIns_3;
  assign io_argIns_2 = regs_io_argIns_4;
  assign io_memStreams_loads_3_cmd_ready = mags_0_io_app_loads_0_cmd_ready;
  assign io_memStreams_loads_3_rdata_valid = mags_0_io_app_loads_0_rdata_valid;
  assign io_memStreams_loads_3_rdata_bits_0 = mags_0_io_app_loads_0_rdata_bits_0;
  assign io_memStreams_loads_2_cmd_ready = mags_1_io_app_loads_0_cmd_ready;
  assign io_memStreams_loads_2_rdata_valid = mags_1_io_app_loads_0_rdata_valid;
  assign io_memStreams_loads_2_rdata_bits_0 = mags_1_io_app_loads_0_rdata_bits_0;
  assign io_memStreams_loads_1_cmd_ready = mags_2_io_app_loads_0_cmd_ready;
  assign io_memStreams_loads_1_rdata_valid = mags_2_io_app_loads_0_rdata_valid;
  assign io_memStreams_loads_1_rdata_bits_0 = mags_2_io_app_loads_0_rdata_bits_0;
  assign io_memStreams_loads_0_cmd_ready = mags_3_io_app_loads_0_cmd_ready;
  assign io_memStreams_loads_0_rdata_valid = mags_3_io_app_loads_0_rdata_valid;
  assign io_memStreams_loads_0_rdata_bits_0 = mags_3_io_app_loads_0_rdata_bits_0;
  assign io_dram_0_cmd_valid = mags_0_io_dram_cmd_valid;
  assign io_dram_0_cmd_bits_addr = mags_0_io_dram_cmd_bits_addr;
  assign io_dram_0_cmd_bits_size = mags_0_io_dram_cmd_bits_size;
  assign io_dram_0_cmd_bits_isWr = mags_0_io_dram_cmd_bits_isWr;
  assign io_dram_0_cmd_bits_tag_uid = mags_0_io_dram_cmd_bits_tag_uid;
  assign io_dram_0_cmd_bits_tag_streamId = mags_0_io_dram_cmd_bits_tag_streamId;
  assign io_dram_0_wdata_valid = mags_0_io_dram_wdata_valid;
  assign io_dram_0_wdata_bits_wdata_0 = mags_0_io_dram_wdata_bits_wdata_0;
  assign io_dram_0_wdata_bits_wdata_1 = mags_0_io_dram_wdata_bits_wdata_1;
  assign io_dram_0_wdata_bits_wdata_2 = mags_0_io_dram_wdata_bits_wdata_2;
  assign io_dram_0_wdata_bits_wdata_3 = mags_0_io_dram_wdata_bits_wdata_3;
  assign io_dram_0_wdata_bits_wdata_4 = mags_0_io_dram_wdata_bits_wdata_4;
  assign io_dram_0_wdata_bits_wdata_5 = mags_0_io_dram_wdata_bits_wdata_5;
  assign io_dram_0_wdata_bits_wdata_6 = mags_0_io_dram_wdata_bits_wdata_6;
  assign io_dram_0_wdata_bits_wdata_7 = mags_0_io_dram_wdata_bits_wdata_7;
  assign io_dram_0_wdata_bits_wdata_8 = mags_0_io_dram_wdata_bits_wdata_8;
  assign io_dram_0_wdata_bits_wdata_9 = mags_0_io_dram_wdata_bits_wdata_9;
  assign io_dram_0_wdata_bits_wdata_10 = mags_0_io_dram_wdata_bits_wdata_10;
  assign io_dram_0_wdata_bits_wdata_11 = mags_0_io_dram_wdata_bits_wdata_11;
  assign io_dram_0_wdata_bits_wdata_12 = mags_0_io_dram_wdata_bits_wdata_12;
  assign io_dram_0_wdata_bits_wdata_13 = mags_0_io_dram_wdata_bits_wdata_13;
  assign io_dram_0_wdata_bits_wdata_14 = mags_0_io_dram_wdata_bits_wdata_14;
  assign io_dram_0_wdata_bits_wdata_15 = mags_0_io_dram_wdata_bits_wdata_15;
  assign io_dram_0_wdata_bits_wstrb_0 = mags_0_io_dram_wdata_bits_wstrb_0;
  assign io_dram_0_wdata_bits_wstrb_1 = mags_0_io_dram_wdata_bits_wstrb_1;
  assign io_dram_0_wdata_bits_wstrb_2 = mags_0_io_dram_wdata_bits_wstrb_2;
  assign io_dram_0_wdata_bits_wstrb_3 = mags_0_io_dram_wdata_bits_wstrb_3;
  assign io_dram_0_wdata_bits_wstrb_4 = mags_0_io_dram_wdata_bits_wstrb_4;
  assign io_dram_0_wdata_bits_wstrb_5 = mags_0_io_dram_wdata_bits_wstrb_5;
  assign io_dram_0_wdata_bits_wstrb_6 = mags_0_io_dram_wdata_bits_wstrb_6;
  assign io_dram_0_wdata_bits_wstrb_7 = mags_0_io_dram_wdata_bits_wstrb_7;
  assign io_dram_0_wdata_bits_wstrb_8 = mags_0_io_dram_wdata_bits_wstrb_8;
  assign io_dram_0_wdata_bits_wstrb_9 = mags_0_io_dram_wdata_bits_wstrb_9;
  assign io_dram_0_wdata_bits_wstrb_10 = mags_0_io_dram_wdata_bits_wstrb_10;
  assign io_dram_0_wdata_bits_wstrb_11 = mags_0_io_dram_wdata_bits_wstrb_11;
  assign io_dram_0_wdata_bits_wstrb_12 = mags_0_io_dram_wdata_bits_wstrb_12;
  assign io_dram_0_wdata_bits_wstrb_13 = mags_0_io_dram_wdata_bits_wstrb_13;
  assign io_dram_0_wdata_bits_wstrb_14 = mags_0_io_dram_wdata_bits_wstrb_14;
  assign io_dram_0_wdata_bits_wstrb_15 = mags_0_io_dram_wdata_bits_wstrb_15;
  assign io_dram_0_wdata_bits_wstrb_16 = mags_0_io_dram_wdata_bits_wstrb_16;
  assign io_dram_0_wdata_bits_wstrb_17 = mags_0_io_dram_wdata_bits_wstrb_17;
  assign io_dram_0_wdata_bits_wstrb_18 = mags_0_io_dram_wdata_bits_wstrb_18;
  assign io_dram_0_wdata_bits_wstrb_19 = mags_0_io_dram_wdata_bits_wstrb_19;
  assign io_dram_0_wdata_bits_wstrb_20 = mags_0_io_dram_wdata_bits_wstrb_20;
  assign io_dram_0_wdata_bits_wstrb_21 = mags_0_io_dram_wdata_bits_wstrb_21;
  assign io_dram_0_wdata_bits_wstrb_22 = mags_0_io_dram_wdata_bits_wstrb_22;
  assign io_dram_0_wdata_bits_wstrb_23 = mags_0_io_dram_wdata_bits_wstrb_23;
  assign io_dram_0_wdata_bits_wstrb_24 = mags_0_io_dram_wdata_bits_wstrb_24;
  assign io_dram_0_wdata_bits_wstrb_25 = mags_0_io_dram_wdata_bits_wstrb_25;
  assign io_dram_0_wdata_bits_wstrb_26 = mags_0_io_dram_wdata_bits_wstrb_26;
  assign io_dram_0_wdata_bits_wstrb_27 = mags_0_io_dram_wdata_bits_wstrb_27;
  assign io_dram_0_wdata_bits_wstrb_28 = mags_0_io_dram_wdata_bits_wstrb_28;
  assign io_dram_0_wdata_bits_wstrb_29 = mags_0_io_dram_wdata_bits_wstrb_29;
  assign io_dram_0_wdata_bits_wstrb_30 = mags_0_io_dram_wdata_bits_wstrb_30;
  assign io_dram_0_wdata_bits_wstrb_31 = mags_0_io_dram_wdata_bits_wstrb_31;
  assign io_dram_0_wdata_bits_wstrb_32 = mags_0_io_dram_wdata_bits_wstrb_32;
  assign io_dram_0_wdata_bits_wstrb_33 = mags_0_io_dram_wdata_bits_wstrb_33;
  assign io_dram_0_wdata_bits_wstrb_34 = mags_0_io_dram_wdata_bits_wstrb_34;
  assign io_dram_0_wdata_bits_wstrb_35 = mags_0_io_dram_wdata_bits_wstrb_35;
  assign io_dram_0_wdata_bits_wstrb_36 = mags_0_io_dram_wdata_bits_wstrb_36;
  assign io_dram_0_wdata_bits_wstrb_37 = mags_0_io_dram_wdata_bits_wstrb_37;
  assign io_dram_0_wdata_bits_wstrb_38 = mags_0_io_dram_wdata_bits_wstrb_38;
  assign io_dram_0_wdata_bits_wstrb_39 = mags_0_io_dram_wdata_bits_wstrb_39;
  assign io_dram_0_wdata_bits_wstrb_40 = mags_0_io_dram_wdata_bits_wstrb_40;
  assign io_dram_0_wdata_bits_wstrb_41 = mags_0_io_dram_wdata_bits_wstrb_41;
  assign io_dram_0_wdata_bits_wstrb_42 = mags_0_io_dram_wdata_bits_wstrb_42;
  assign io_dram_0_wdata_bits_wstrb_43 = mags_0_io_dram_wdata_bits_wstrb_43;
  assign io_dram_0_wdata_bits_wstrb_44 = mags_0_io_dram_wdata_bits_wstrb_44;
  assign io_dram_0_wdata_bits_wstrb_45 = mags_0_io_dram_wdata_bits_wstrb_45;
  assign io_dram_0_wdata_bits_wstrb_46 = mags_0_io_dram_wdata_bits_wstrb_46;
  assign io_dram_0_wdata_bits_wstrb_47 = mags_0_io_dram_wdata_bits_wstrb_47;
  assign io_dram_0_wdata_bits_wstrb_48 = mags_0_io_dram_wdata_bits_wstrb_48;
  assign io_dram_0_wdata_bits_wstrb_49 = mags_0_io_dram_wdata_bits_wstrb_49;
  assign io_dram_0_wdata_bits_wstrb_50 = mags_0_io_dram_wdata_bits_wstrb_50;
  assign io_dram_0_wdata_bits_wstrb_51 = mags_0_io_dram_wdata_bits_wstrb_51;
  assign io_dram_0_wdata_bits_wstrb_52 = mags_0_io_dram_wdata_bits_wstrb_52;
  assign io_dram_0_wdata_bits_wstrb_53 = mags_0_io_dram_wdata_bits_wstrb_53;
  assign io_dram_0_wdata_bits_wstrb_54 = mags_0_io_dram_wdata_bits_wstrb_54;
  assign io_dram_0_wdata_bits_wstrb_55 = mags_0_io_dram_wdata_bits_wstrb_55;
  assign io_dram_0_wdata_bits_wstrb_56 = mags_0_io_dram_wdata_bits_wstrb_56;
  assign io_dram_0_wdata_bits_wstrb_57 = mags_0_io_dram_wdata_bits_wstrb_57;
  assign io_dram_0_wdata_bits_wstrb_58 = mags_0_io_dram_wdata_bits_wstrb_58;
  assign io_dram_0_wdata_bits_wstrb_59 = mags_0_io_dram_wdata_bits_wstrb_59;
  assign io_dram_0_wdata_bits_wstrb_60 = mags_0_io_dram_wdata_bits_wstrb_60;
  assign io_dram_0_wdata_bits_wstrb_61 = mags_0_io_dram_wdata_bits_wstrb_61;
  assign io_dram_0_wdata_bits_wstrb_62 = mags_0_io_dram_wdata_bits_wstrb_62;
  assign io_dram_0_wdata_bits_wstrb_63 = mags_0_io_dram_wdata_bits_wstrb_63;
  assign io_dram_0_rresp_ready = mags_0_io_dram_rresp_ready;
  assign io_dram_0_wresp_ready = mags_0_io_dram_wresp_ready;
  assign io_dram_1_cmd_valid = mags_1_io_dram_cmd_valid;
  assign io_dram_1_cmd_bits_addr = mags_1_io_dram_cmd_bits_addr;
  assign io_dram_1_cmd_bits_size = mags_1_io_dram_cmd_bits_size;
  assign io_dram_1_cmd_bits_isWr = mags_1_io_dram_cmd_bits_isWr;
  assign io_dram_1_cmd_bits_tag_uid = mags_1_io_dram_cmd_bits_tag_uid;
  assign io_dram_1_cmd_bits_tag_streamId = mags_1_io_dram_cmd_bits_tag_streamId;
  assign io_dram_1_wdata_valid = mags_1_io_dram_wdata_valid;
  assign io_dram_1_wdata_bits_wdata_0 = mags_1_io_dram_wdata_bits_wdata_0;
  assign io_dram_1_wdata_bits_wdata_1 = mags_1_io_dram_wdata_bits_wdata_1;
  assign io_dram_1_wdata_bits_wdata_2 = mags_1_io_dram_wdata_bits_wdata_2;
  assign io_dram_1_wdata_bits_wdata_3 = mags_1_io_dram_wdata_bits_wdata_3;
  assign io_dram_1_wdata_bits_wdata_4 = mags_1_io_dram_wdata_bits_wdata_4;
  assign io_dram_1_wdata_bits_wdata_5 = mags_1_io_dram_wdata_bits_wdata_5;
  assign io_dram_1_wdata_bits_wdata_6 = mags_1_io_dram_wdata_bits_wdata_6;
  assign io_dram_1_wdata_bits_wdata_7 = mags_1_io_dram_wdata_bits_wdata_7;
  assign io_dram_1_wdata_bits_wdata_8 = mags_1_io_dram_wdata_bits_wdata_8;
  assign io_dram_1_wdata_bits_wdata_9 = mags_1_io_dram_wdata_bits_wdata_9;
  assign io_dram_1_wdata_bits_wdata_10 = mags_1_io_dram_wdata_bits_wdata_10;
  assign io_dram_1_wdata_bits_wdata_11 = mags_1_io_dram_wdata_bits_wdata_11;
  assign io_dram_1_wdata_bits_wdata_12 = mags_1_io_dram_wdata_bits_wdata_12;
  assign io_dram_1_wdata_bits_wdata_13 = mags_1_io_dram_wdata_bits_wdata_13;
  assign io_dram_1_wdata_bits_wdata_14 = mags_1_io_dram_wdata_bits_wdata_14;
  assign io_dram_1_wdata_bits_wdata_15 = mags_1_io_dram_wdata_bits_wdata_15;
  assign io_dram_1_wdata_bits_wstrb_0 = mags_1_io_dram_wdata_bits_wstrb_0;
  assign io_dram_1_wdata_bits_wstrb_1 = mags_1_io_dram_wdata_bits_wstrb_1;
  assign io_dram_1_wdata_bits_wstrb_2 = mags_1_io_dram_wdata_bits_wstrb_2;
  assign io_dram_1_wdata_bits_wstrb_3 = mags_1_io_dram_wdata_bits_wstrb_3;
  assign io_dram_1_wdata_bits_wstrb_4 = mags_1_io_dram_wdata_bits_wstrb_4;
  assign io_dram_1_wdata_bits_wstrb_5 = mags_1_io_dram_wdata_bits_wstrb_5;
  assign io_dram_1_wdata_bits_wstrb_6 = mags_1_io_dram_wdata_bits_wstrb_6;
  assign io_dram_1_wdata_bits_wstrb_7 = mags_1_io_dram_wdata_bits_wstrb_7;
  assign io_dram_1_wdata_bits_wstrb_8 = mags_1_io_dram_wdata_bits_wstrb_8;
  assign io_dram_1_wdata_bits_wstrb_9 = mags_1_io_dram_wdata_bits_wstrb_9;
  assign io_dram_1_wdata_bits_wstrb_10 = mags_1_io_dram_wdata_bits_wstrb_10;
  assign io_dram_1_wdata_bits_wstrb_11 = mags_1_io_dram_wdata_bits_wstrb_11;
  assign io_dram_1_wdata_bits_wstrb_12 = mags_1_io_dram_wdata_bits_wstrb_12;
  assign io_dram_1_wdata_bits_wstrb_13 = mags_1_io_dram_wdata_bits_wstrb_13;
  assign io_dram_1_wdata_bits_wstrb_14 = mags_1_io_dram_wdata_bits_wstrb_14;
  assign io_dram_1_wdata_bits_wstrb_15 = mags_1_io_dram_wdata_bits_wstrb_15;
  assign io_dram_1_wdata_bits_wstrb_16 = mags_1_io_dram_wdata_bits_wstrb_16;
  assign io_dram_1_wdata_bits_wstrb_17 = mags_1_io_dram_wdata_bits_wstrb_17;
  assign io_dram_1_wdata_bits_wstrb_18 = mags_1_io_dram_wdata_bits_wstrb_18;
  assign io_dram_1_wdata_bits_wstrb_19 = mags_1_io_dram_wdata_bits_wstrb_19;
  assign io_dram_1_wdata_bits_wstrb_20 = mags_1_io_dram_wdata_bits_wstrb_20;
  assign io_dram_1_wdata_bits_wstrb_21 = mags_1_io_dram_wdata_bits_wstrb_21;
  assign io_dram_1_wdata_bits_wstrb_22 = mags_1_io_dram_wdata_bits_wstrb_22;
  assign io_dram_1_wdata_bits_wstrb_23 = mags_1_io_dram_wdata_bits_wstrb_23;
  assign io_dram_1_wdata_bits_wstrb_24 = mags_1_io_dram_wdata_bits_wstrb_24;
  assign io_dram_1_wdata_bits_wstrb_25 = mags_1_io_dram_wdata_bits_wstrb_25;
  assign io_dram_1_wdata_bits_wstrb_26 = mags_1_io_dram_wdata_bits_wstrb_26;
  assign io_dram_1_wdata_bits_wstrb_27 = mags_1_io_dram_wdata_bits_wstrb_27;
  assign io_dram_1_wdata_bits_wstrb_28 = mags_1_io_dram_wdata_bits_wstrb_28;
  assign io_dram_1_wdata_bits_wstrb_29 = mags_1_io_dram_wdata_bits_wstrb_29;
  assign io_dram_1_wdata_bits_wstrb_30 = mags_1_io_dram_wdata_bits_wstrb_30;
  assign io_dram_1_wdata_bits_wstrb_31 = mags_1_io_dram_wdata_bits_wstrb_31;
  assign io_dram_1_wdata_bits_wstrb_32 = mags_1_io_dram_wdata_bits_wstrb_32;
  assign io_dram_1_wdata_bits_wstrb_33 = mags_1_io_dram_wdata_bits_wstrb_33;
  assign io_dram_1_wdata_bits_wstrb_34 = mags_1_io_dram_wdata_bits_wstrb_34;
  assign io_dram_1_wdata_bits_wstrb_35 = mags_1_io_dram_wdata_bits_wstrb_35;
  assign io_dram_1_wdata_bits_wstrb_36 = mags_1_io_dram_wdata_bits_wstrb_36;
  assign io_dram_1_wdata_bits_wstrb_37 = mags_1_io_dram_wdata_bits_wstrb_37;
  assign io_dram_1_wdata_bits_wstrb_38 = mags_1_io_dram_wdata_bits_wstrb_38;
  assign io_dram_1_wdata_bits_wstrb_39 = mags_1_io_dram_wdata_bits_wstrb_39;
  assign io_dram_1_wdata_bits_wstrb_40 = mags_1_io_dram_wdata_bits_wstrb_40;
  assign io_dram_1_wdata_bits_wstrb_41 = mags_1_io_dram_wdata_bits_wstrb_41;
  assign io_dram_1_wdata_bits_wstrb_42 = mags_1_io_dram_wdata_bits_wstrb_42;
  assign io_dram_1_wdata_bits_wstrb_43 = mags_1_io_dram_wdata_bits_wstrb_43;
  assign io_dram_1_wdata_bits_wstrb_44 = mags_1_io_dram_wdata_bits_wstrb_44;
  assign io_dram_1_wdata_bits_wstrb_45 = mags_1_io_dram_wdata_bits_wstrb_45;
  assign io_dram_1_wdata_bits_wstrb_46 = mags_1_io_dram_wdata_bits_wstrb_46;
  assign io_dram_1_wdata_bits_wstrb_47 = mags_1_io_dram_wdata_bits_wstrb_47;
  assign io_dram_1_wdata_bits_wstrb_48 = mags_1_io_dram_wdata_bits_wstrb_48;
  assign io_dram_1_wdata_bits_wstrb_49 = mags_1_io_dram_wdata_bits_wstrb_49;
  assign io_dram_1_wdata_bits_wstrb_50 = mags_1_io_dram_wdata_bits_wstrb_50;
  assign io_dram_1_wdata_bits_wstrb_51 = mags_1_io_dram_wdata_bits_wstrb_51;
  assign io_dram_1_wdata_bits_wstrb_52 = mags_1_io_dram_wdata_bits_wstrb_52;
  assign io_dram_1_wdata_bits_wstrb_53 = mags_1_io_dram_wdata_bits_wstrb_53;
  assign io_dram_1_wdata_bits_wstrb_54 = mags_1_io_dram_wdata_bits_wstrb_54;
  assign io_dram_1_wdata_bits_wstrb_55 = mags_1_io_dram_wdata_bits_wstrb_55;
  assign io_dram_1_wdata_bits_wstrb_56 = mags_1_io_dram_wdata_bits_wstrb_56;
  assign io_dram_1_wdata_bits_wstrb_57 = mags_1_io_dram_wdata_bits_wstrb_57;
  assign io_dram_1_wdata_bits_wstrb_58 = mags_1_io_dram_wdata_bits_wstrb_58;
  assign io_dram_1_wdata_bits_wstrb_59 = mags_1_io_dram_wdata_bits_wstrb_59;
  assign io_dram_1_wdata_bits_wstrb_60 = mags_1_io_dram_wdata_bits_wstrb_60;
  assign io_dram_1_wdata_bits_wstrb_61 = mags_1_io_dram_wdata_bits_wstrb_61;
  assign io_dram_1_wdata_bits_wstrb_62 = mags_1_io_dram_wdata_bits_wstrb_62;
  assign io_dram_1_wdata_bits_wstrb_63 = mags_1_io_dram_wdata_bits_wstrb_63;
  assign io_dram_1_rresp_ready = mags_1_io_dram_rresp_ready;
  assign io_dram_1_wresp_ready = mags_1_io_dram_wresp_ready;
  assign io_dram_2_cmd_valid = mags_2_io_dram_cmd_valid;
  assign io_dram_2_cmd_bits_addr = mags_2_io_dram_cmd_bits_addr;
  assign io_dram_2_cmd_bits_size = mags_2_io_dram_cmd_bits_size;
  assign io_dram_2_cmd_bits_isWr = mags_2_io_dram_cmd_bits_isWr;
  assign io_dram_2_cmd_bits_tag_uid = mags_2_io_dram_cmd_bits_tag_uid;
  assign io_dram_2_cmd_bits_tag_streamId = mags_2_io_dram_cmd_bits_tag_streamId;
  assign io_dram_2_wdata_valid = mags_2_io_dram_wdata_valid;
  assign io_dram_2_wdata_bits_wdata_0 = mags_2_io_dram_wdata_bits_wdata_0;
  assign io_dram_2_wdata_bits_wdata_1 = mags_2_io_dram_wdata_bits_wdata_1;
  assign io_dram_2_wdata_bits_wdata_2 = mags_2_io_dram_wdata_bits_wdata_2;
  assign io_dram_2_wdata_bits_wdata_3 = mags_2_io_dram_wdata_bits_wdata_3;
  assign io_dram_2_wdata_bits_wdata_4 = mags_2_io_dram_wdata_bits_wdata_4;
  assign io_dram_2_wdata_bits_wdata_5 = mags_2_io_dram_wdata_bits_wdata_5;
  assign io_dram_2_wdata_bits_wdata_6 = mags_2_io_dram_wdata_bits_wdata_6;
  assign io_dram_2_wdata_bits_wdata_7 = mags_2_io_dram_wdata_bits_wdata_7;
  assign io_dram_2_wdata_bits_wdata_8 = mags_2_io_dram_wdata_bits_wdata_8;
  assign io_dram_2_wdata_bits_wdata_9 = mags_2_io_dram_wdata_bits_wdata_9;
  assign io_dram_2_wdata_bits_wdata_10 = mags_2_io_dram_wdata_bits_wdata_10;
  assign io_dram_2_wdata_bits_wdata_11 = mags_2_io_dram_wdata_bits_wdata_11;
  assign io_dram_2_wdata_bits_wdata_12 = mags_2_io_dram_wdata_bits_wdata_12;
  assign io_dram_2_wdata_bits_wdata_13 = mags_2_io_dram_wdata_bits_wdata_13;
  assign io_dram_2_wdata_bits_wdata_14 = mags_2_io_dram_wdata_bits_wdata_14;
  assign io_dram_2_wdata_bits_wdata_15 = mags_2_io_dram_wdata_bits_wdata_15;
  assign io_dram_2_wdata_bits_wstrb_0 = mags_2_io_dram_wdata_bits_wstrb_0;
  assign io_dram_2_wdata_bits_wstrb_1 = mags_2_io_dram_wdata_bits_wstrb_1;
  assign io_dram_2_wdata_bits_wstrb_2 = mags_2_io_dram_wdata_bits_wstrb_2;
  assign io_dram_2_wdata_bits_wstrb_3 = mags_2_io_dram_wdata_bits_wstrb_3;
  assign io_dram_2_wdata_bits_wstrb_4 = mags_2_io_dram_wdata_bits_wstrb_4;
  assign io_dram_2_wdata_bits_wstrb_5 = mags_2_io_dram_wdata_bits_wstrb_5;
  assign io_dram_2_wdata_bits_wstrb_6 = mags_2_io_dram_wdata_bits_wstrb_6;
  assign io_dram_2_wdata_bits_wstrb_7 = mags_2_io_dram_wdata_bits_wstrb_7;
  assign io_dram_2_wdata_bits_wstrb_8 = mags_2_io_dram_wdata_bits_wstrb_8;
  assign io_dram_2_wdata_bits_wstrb_9 = mags_2_io_dram_wdata_bits_wstrb_9;
  assign io_dram_2_wdata_bits_wstrb_10 = mags_2_io_dram_wdata_bits_wstrb_10;
  assign io_dram_2_wdata_bits_wstrb_11 = mags_2_io_dram_wdata_bits_wstrb_11;
  assign io_dram_2_wdata_bits_wstrb_12 = mags_2_io_dram_wdata_bits_wstrb_12;
  assign io_dram_2_wdata_bits_wstrb_13 = mags_2_io_dram_wdata_bits_wstrb_13;
  assign io_dram_2_wdata_bits_wstrb_14 = mags_2_io_dram_wdata_bits_wstrb_14;
  assign io_dram_2_wdata_bits_wstrb_15 = mags_2_io_dram_wdata_bits_wstrb_15;
  assign io_dram_2_wdata_bits_wstrb_16 = mags_2_io_dram_wdata_bits_wstrb_16;
  assign io_dram_2_wdata_bits_wstrb_17 = mags_2_io_dram_wdata_bits_wstrb_17;
  assign io_dram_2_wdata_bits_wstrb_18 = mags_2_io_dram_wdata_bits_wstrb_18;
  assign io_dram_2_wdata_bits_wstrb_19 = mags_2_io_dram_wdata_bits_wstrb_19;
  assign io_dram_2_wdata_bits_wstrb_20 = mags_2_io_dram_wdata_bits_wstrb_20;
  assign io_dram_2_wdata_bits_wstrb_21 = mags_2_io_dram_wdata_bits_wstrb_21;
  assign io_dram_2_wdata_bits_wstrb_22 = mags_2_io_dram_wdata_bits_wstrb_22;
  assign io_dram_2_wdata_bits_wstrb_23 = mags_2_io_dram_wdata_bits_wstrb_23;
  assign io_dram_2_wdata_bits_wstrb_24 = mags_2_io_dram_wdata_bits_wstrb_24;
  assign io_dram_2_wdata_bits_wstrb_25 = mags_2_io_dram_wdata_bits_wstrb_25;
  assign io_dram_2_wdata_bits_wstrb_26 = mags_2_io_dram_wdata_bits_wstrb_26;
  assign io_dram_2_wdata_bits_wstrb_27 = mags_2_io_dram_wdata_bits_wstrb_27;
  assign io_dram_2_wdata_bits_wstrb_28 = mags_2_io_dram_wdata_bits_wstrb_28;
  assign io_dram_2_wdata_bits_wstrb_29 = mags_2_io_dram_wdata_bits_wstrb_29;
  assign io_dram_2_wdata_bits_wstrb_30 = mags_2_io_dram_wdata_bits_wstrb_30;
  assign io_dram_2_wdata_bits_wstrb_31 = mags_2_io_dram_wdata_bits_wstrb_31;
  assign io_dram_2_wdata_bits_wstrb_32 = mags_2_io_dram_wdata_bits_wstrb_32;
  assign io_dram_2_wdata_bits_wstrb_33 = mags_2_io_dram_wdata_bits_wstrb_33;
  assign io_dram_2_wdata_bits_wstrb_34 = mags_2_io_dram_wdata_bits_wstrb_34;
  assign io_dram_2_wdata_bits_wstrb_35 = mags_2_io_dram_wdata_bits_wstrb_35;
  assign io_dram_2_wdata_bits_wstrb_36 = mags_2_io_dram_wdata_bits_wstrb_36;
  assign io_dram_2_wdata_bits_wstrb_37 = mags_2_io_dram_wdata_bits_wstrb_37;
  assign io_dram_2_wdata_bits_wstrb_38 = mags_2_io_dram_wdata_bits_wstrb_38;
  assign io_dram_2_wdata_bits_wstrb_39 = mags_2_io_dram_wdata_bits_wstrb_39;
  assign io_dram_2_wdata_bits_wstrb_40 = mags_2_io_dram_wdata_bits_wstrb_40;
  assign io_dram_2_wdata_bits_wstrb_41 = mags_2_io_dram_wdata_bits_wstrb_41;
  assign io_dram_2_wdata_bits_wstrb_42 = mags_2_io_dram_wdata_bits_wstrb_42;
  assign io_dram_2_wdata_bits_wstrb_43 = mags_2_io_dram_wdata_bits_wstrb_43;
  assign io_dram_2_wdata_bits_wstrb_44 = mags_2_io_dram_wdata_bits_wstrb_44;
  assign io_dram_2_wdata_bits_wstrb_45 = mags_2_io_dram_wdata_bits_wstrb_45;
  assign io_dram_2_wdata_bits_wstrb_46 = mags_2_io_dram_wdata_bits_wstrb_46;
  assign io_dram_2_wdata_bits_wstrb_47 = mags_2_io_dram_wdata_bits_wstrb_47;
  assign io_dram_2_wdata_bits_wstrb_48 = mags_2_io_dram_wdata_bits_wstrb_48;
  assign io_dram_2_wdata_bits_wstrb_49 = mags_2_io_dram_wdata_bits_wstrb_49;
  assign io_dram_2_wdata_bits_wstrb_50 = mags_2_io_dram_wdata_bits_wstrb_50;
  assign io_dram_2_wdata_bits_wstrb_51 = mags_2_io_dram_wdata_bits_wstrb_51;
  assign io_dram_2_wdata_bits_wstrb_52 = mags_2_io_dram_wdata_bits_wstrb_52;
  assign io_dram_2_wdata_bits_wstrb_53 = mags_2_io_dram_wdata_bits_wstrb_53;
  assign io_dram_2_wdata_bits_wstrb_54 = mags_2_io_dram_wdata_bits_wstrb_54;
  assign io_dram_2_wdata_bits_wstrb_55 = mags_2_io_dram_wdata_bits_wstrb_55;
  assign io_dram_2_wdata_bits_wstrb_56 = mags_2_io_dram_wdata_bits_wstrb_56;
  assign io_dram_2_wdata_bits_wstrb_57 = mags_2_io_dram_wdata_bits_wstrb_57;
  assign io_dram_2_wdata_bits_wstrb_58 = mags_2_io_dram_wdata_bits_wstrb_58;
  assign io_dram_2_wdata_bits_wstrb_59 = mags_2_io_dram_wdata_bits_wstrb_59;
  assign io_dram_2_wdata_bits_wstrb_60 = mags_2_io_dram_wdata_bits_wstrb_60;
  assign io_dram_2_wdata_bits_wstrb_61 = mags_2_io_dram_wdata_bits_wstrb_61;
  assign io_dram_2_wdata_bits_wstrb_62 = mags_2_io_dram_wdata_bits_wstrb_62;
  assign io_dram_2_wdata_bits_wstrb_63 = mags_2_io_dram_wdata_bits_wstrb_63;
  assign io_dram_2_rresp_ready = mags_2_io_dram_rresp_ready;
  assign io_dram_2_wresp_ready = mags_2_io_dram_wresp_ready;
  assign io_dram_3_cmd_valid = mags_3_io_dram_cmd_valid;
  assign io_dram_3_cmd_bits_addr = mags_3_io_dram_cmd_bits_addr;
  assign io_dram_3_cmd_bits_size = mags_3_io_dram_cmd_bits_size;
  assign io_dram_3_cmd_bits_isWr = mags_3_io_dram_cmd_bits_isWr;
  assign io_dram_3_cmd_bits_tag_uid = mags_3_io_dram_cmd_bits_tag_uid;
  assign io_dram_3_cmd_bits_tag_streamId = mags_3_io_dram_cmd_bits_tag_streamId;
  assign io_dram_3_wdata_valid = mags_3_io_dram_wdata_valid;
  assign io_dram_3_wdata_bits_wdata_0 = mags_3_io_dram_wdata_bits_wdata_0;
  assign io_dram_3_wdata_bits_wdata_1 = mags_3_io_dram_wdata_bits_wdata_1;
  assign io_dram_3_wdata_bits_wdata_2 = mags_3_io_dram_wdata_bits_wdata_2;
  assign io_dram_3_wdata_bits_wdata_3 = mags_3_io_dram_wdata_bits_wdata_3;
  assign io_dram_3_wdata_bits_wdata_4 = mags_3_io_dram_wdata_bits_wdata_4;
  assign io_dram_3_wdata_bits_wdata_5 = mags_3_io_dram_wdata_bits_wdata_5;
  assign io_dram_3_wdata_bits_wdata_6 = mags_3_io_dram_wdata_bits_wdata_6;
  assign io_dram_3_wdata_bits_wdata_7 = mags_3_io_dram_wdata_bits_wdata_7;
  assign io_dram_3_wdata_bits_wdata_8 = mags_3_io_dram_wdata_bits_wdata_8;
  assign io_dram_3_wdata_bits_wdata_9 = mags_3_io_dram_wdata_bits_wdata_9;
  assign io_dram_3_wdata_bits_wdata_10 = mags_3_io_dram_wdata_bits_wdata_10;
  assign io_dram_3_wdata_bits_wdata_11 = mags_3_io_dram_wdata_bits_wdata_11;
  assign io_dram_3_wdata_bits_wdata_12 = mags_3_io_dram_wdata_bits_wdata_12;
  assign io_dram_3_wdata_bits_wdata_13 = mags_3_io_dram_wdata_bits_wdata_13;
  assign io_dram_3_wdata_bits_wdata_14 = mags_3_io_dram_wdata_bits_wdata_14;
  assign io_dram_3_wdata_bits_wdata_15 = mags_3_io_dram_wdata_bits_wdata_15;
  assign io_dram_3_wdata_bits_wstrb_0 = mags_3_io_dram_wdata_bits_wstrb_0;
  assign io_dram_3_wdata_bits_wstrb_1 = mags_3_io_dram_wdata_bits_wstrb_1;
  assign io_dram_3_wdata_bits_wstrb_2 = mags_3_io_dram_wdata_bits_wstrb_2;
  assign io_dram_3_wdata_bits_wstrb_3 = mags_3_io_dram_wdata_bits_wstrb_3;
  assign io_dram_3_wdata_bits_wstrb_4 = mags_3_io_dram_wdata_bits_wstrb_4;
  assign io_dram_3_wdata_bits_wstrb_5 = mags_3_io_dram_wdata_bits_wstrb_5;
  assign io_dram_3_wdata_bits_wstrb_6 = mags_3_io_dram_wdata_bits_wstrb_6;
  assign io_dram_3_wdata_bits_wstrb_7 = mags_3_io_dram_wdata_bits_wstrb_7;
  assign io_dram_3_wdata_bits_wstrb_8 = mags_3_io_dram_wdata_bits_wstrb_8;
  assign io_dram_3_wdata_bits_wstrb_9 = mags_3_io_dram_wdata_bits_wstrb_9;
  assign io_dram_3_wdata_bits_wstrb_10 = mags_3_io_dram_wdata_bits_wstrb_10;
  assign io_dram_3_wdata_bits_wstrb_11 = mags_3_io_dram_wdata_bits_wstrb_11;
  assign io_dram_3_wdata_bits_wstrb_12 = mags_3_io_dram_wdata_bits_wstrb_12;
  assign io_dram_3_wdata_bits_wstrb_13 = mags_3_io_dram_wdata_bits_wstrb_13;
  assign io_dram_3_wdata_bits_wstrb_14 = mags_3_io_dram_wdata_bits_wstrb_14;
  assign io_dram_3_wdata_bits_wstrb_15 = mags_3_io_dram_wdata_bits_wstrb_15;
  assign io_dram_3_wdata_bits_wstrb_16 = mags_3_io_dram_wdata_bits_wstrb_16;
  assign io_dram_3_wdata_bits_wstrb_17 = mags_3_io_dram_wdata_bits_wstrb_17;
  assign io_dram_3_wdata_bits_wstrb_18 = mags_3_io_dram_wdata_bits_wstrb_18;
  assign io_dram_3_wdata_bits_wstrb_19 = mags_3_io_dram_wdata_bits_wstrb_19;
  assign io_dram_3_wdata_bits_wstrb_20 = mags_3_io_dram_wdata_bits_wstrb_20;
  assign io_dram_3_wdata_bits_wstrb_21 = mags_3_io_dram_wdata_bits_wstrb_21;
  assign io_dram_3_wdata_bits_wstrb_22 = mags_3_io_dram_wdata_bits_wstrb_22;
  assign io_dram_3_wdata_bits_wstrb_23 = mags_3_io_dram_wdata_bits_wstrb_23;
  assign io_dram_3_wdata_bits_wstrb_24 = mags_3_io_dram_wdata_bits_wstrb_24;
  assign io_dram_3_wdata_bits_wstrb_25 = mags_3_io_dram_wdata_bits_wstrb_25;
  assign io_dram_3_wdata_bits_wstrb_26 = mags_3_io_dram_wdata_bits_wstrb_26;
  assign io_dram_3_wdata_bits_wstrb_27 = mags_3_io_dram_wdata_bits_wstrb_27;
  assign io_dram_3_wdata_bits_wstrb_28 = mags_3_io_dram_wdata_bits_wstrb_28;
  assign io_dram_3_wdata_bits_wstrb_29 = mags_3_io_dram_wdata_bits_wstrb_29;
  assign io_dram_3_wdata_bits_wstrb_30 = mags_3_io_dram_wdata_bits_wstrb_30;
  assign io_dram_3_wdata_bits_wstrb_31 = mags_3_io_dram_wdata_bits_wstrb_31;
  assign io_dram_3_wdata_bits_wstrb_32 = mags_3_io_dram_wdata_bits_wstrb_32;
  assign io_dram_3_wdata_bits_wstrb_33 = mags_3_io_dram_wdata_bits_wstrb_33;
  assign io_dram_3_wdata_bits_wstrb_34 = mags_3_io_dram_wdata_bits_wstrb_34;
  assign io_dram_3_wdata_bits_wstrb_35 = mags_3_io_dram_wdata_bits_wstrb_35;
  assign io_dram_3_wdata_bits_wstrb_36 = mags_3_io_dram_wdata_bits_wstrb_36;
  assign io_dram_3_wdata_bits_wstrb_37 = mags_3_io_dram_wdata_bits_wstrb_37;
  assign io_dram_3_wdata_bits_wstrb_38 = mags_3_io_dram_wdata_bits_wstrb_38;
  assign io_dram_3_wdata_bits_wstrb_39 = mags_3_io_dram_wdata_bits_wstrb_39;
  assign io_dram_3_wdata_bits_wstrb_40 = mags_3_io_dram_wdata_bits_wstrb_40;
  assign io_dram_3_wdata_bits_wstrb_41 = mags_3_io_dram_wdata_bits_wstrb_41;
  assign io_dram_3_wdata_bits_wstrb_42 = mags_3_io_dram_wdata_bits_wstrb_42;
  assign io_dram_3_wdata_bits_wstrb_43 = mags_3_io_dram_wdata_bits_wstrb_43;
  assign io_dram_3_wdata_bits_wstrb_44 = mags_3_io_dram_wdata_bits_wstrb_44;
  assign io_dram_3_wdata_bits_wstrb_45 = mags_3_io_dram_wdata_bits_wstrb_45;
  assign io_dram_3_wdata_bits_wstrb_46 = mags_3_io_dram_wdata_bits_wstrb_46;
  assign io_dram_3_wdata_bits_wstrb_47 = mags_3_io_dram_wdata_bits_wstrb_47;
  assign io_dram_3_wdata_bits_wstrb_48 = mags_3_io_dram_wdata_bits_wstrb_48;
  assign io_dram_3_wdata_bits_wstrb_49 = mags_3_io_dram_wdata_bits_wstrb_49;
  assign io_dram_3_wdata_bits_wstrb_50 = mags_3_io_dram_wdata_bits_wstrb_50;
  assign io_dram_3_wdata_bits_wstrb_51 = mags_3_io_dram_wdata_bits_wstrb_51;
  assign io_dram_3_wdata_bits_wstrb_52 = mags_3_io_dram_wdata_bits_wstrb_52;
  assign io_dram_3_wdata_bits_wstrb_53 = mags_3_io_dram_wdata_bits_wstrb_53;
  assign io_dram_3_wdata_bits_wstrb_54 = mags_3_io_dram_wdata_bits_wstrb_54;
  assign io_dram_3_wdata_bits_wstrb_55 = mags_3_io_dram_wdata_bits_wstrb_55;
  assign io_dram_3_wdata_bits_wstrb_56 = mags_3_io_dram_wdata_bits_wstrb_56;
  assign io_dram_3_wdata_bits_wstrb_57 = mags_3_io_dram_wdata_bits_wstrb_57;
  assign io_dram_3_wdata_bits_wstrb_58 = mags_3_io_dram_wdata_bits_wstrb_58;
  assign io_dram_3_wdata_bits_wstrb_59 = mags_3_io_dram_wdata_bits_wstrb_59;
  assign io_dram_3_wdata_bits_wstrb_60 = mags_3_io_dram_wdata_bits_wstrb_60;
  assign io_dram_3_wdata_bits_wstrb_61 = mags_3_io_dram_wdata_bits_wstrb_61;
  assign io_dram_3_wdata_bits_wstrb_62 = mags_3_io_dram_wdata_bits_wstrb_62;
  assign io_dram_3_wdata_bits_wstrb_63 = mags_3_io_dram_wdata_bits_wstrb_63;
  assign io_dram_3_rresp_ready = mags_3_io_dram_rresp_ready;
  assign io_dram_3_wresp_ready = mags_3_io_dram_wresp_ready;
  assign mags_0_io_enable = localEnable;
  assign mags_0_io_reset = localReset;
  assign mags_0_io_app_loads_0_cmd_valid = io_memStreams_loads_3_cmd_valid;
  assign mags_0_io_app_loads_0_cmd_bits_addr = io_memStreams_loads_3_cmd_bits_addr;
  assign mags_0_io_app_loads_0_cmd_bits_isWr = io_memStreams_loads_3_cmd_bits_isWr;
  assign mags_0_io_app_loads_0_cmd_bits_size = io_memStreams_loads_3_cmd_bits_size;
  assign mags_0_io_app_loads_0_rdata_ready = io_memStreams_loads_3_rdata_ready;
  assign mags_0_io_dram_cmd_ready = io_dram_0_cmd_ready;
  assign mags_0_io_dram_wdata_ready = io_dram_0_wdata_ready;
  assign mags_0_io_dram_rresp_valid = io_dram_0_rresp_valid;
  assign mags_0_io_dram_rresp_bits_rdata_0 = io_dram_0_rresp_bits_rdata_0;
  assign mags_0_io_dram_rresp_bits_rdata_1 = io_dram_0_rresp_bits_rdata_1;
  assign mags_0_io_dram_rresp_bits_rdata_2 = io_dram_0_rresp_bits_rdata_2;
  assign mags_0_io_dram_rresp_bits_rdata_3 = io_dram_0_rresp_bits_rdata_3;
  assign mags_0_io_dram_rresp_bits_rdata_4 = io_dram_0_rresp_bits_rdata_4;
  assign mags_0_io_dram_rresp_bits_rdata_5 = io_dram_0_rresp_bits_rdata_5;
  assign mags_0_io_dram_rresp_bits_rdata_6 = io_dram_0_rresp_bits_rdata_6;
  assign mags_0_io_dram_rresp_bits_rdata_7 = io_dram_0_rresp_bits_rdata_7;
  assign mags_0_io_dram_rresp_bits_rdata_8 = io_dram_0_rresp_bits_rdata_8;
  assign mags_0_io_dram_rresp_bits_rdata_9 = io_dram_0_rresp_bits_rdata_9;
  assign mags_0_io_dram_rresp_bits_rdata_10 = io_dram_0_rresp_bits_rdata_10;
  assign mags_0_io_dram_rresp_bits_rdata_11 = io_dram_0_rresp_bits_rdata_11;
  assign mags_0_io_dram_rresp_bits_rdata_12 = io_dram_0_rresp_bits_rdata_12;
  assign mags_0_io_dram_rresp_bits_rdata_13 = io_dram_0_rresp_bits_rdata_13;
  assign mags_0_io_dram_rresp_bits_rdata_14 = io_dram_0_rresp_bits_rdata_14;
  assign mags_0_io_dram_rresp_bits_rdata_15 = io_dram_0_rresp_bits_rdata_15;
  assign mags_0_io_dram_rresp_bits_tag_streamId = io_dram_0_rresp_bits_tag_streamId;
  assign mags_0_io_dram_wresp_valid = io_dram_0_wresp_valid;
  assign mags_0_io_dram_wresp_bits_tag_streamId = io_dram_0_wresp_bits_tag_streamId;
  assign mags_0_io_TOP_AXI_AWADDR = io_TOP_AXI_AWADDR;
  assign mags_0_io_TOP_AXI_AWLEN = io_TOP_AXI_AWLEN;
  assign mags_0_io_TOP_AXI_AWVALID = io_TOP_AXI_AWVALID;
  assign mags_0_io_TOP_AXI_AWREADY = io_TOP_AXI_AWREADY;
  assign mags_0_io_TOP_AXI_ARID = io_TOP_AXI_ARID;
  assign mags_0_io_TOP_AXI_ARADDR = io_TOP_AXI_ARADDR;
  assign mags_0_io_TOP_AXI_ARLEN = io_TOP_AXI_ARLEN;
  assign mags_0_io_TOP_AXI_ARSIZE = io_TOP_AXI_ARSIZE;
  assign mags_0_io_TOP_AXI_ARBURST = io_TOP_AXI_ARBURST;
  assign mags_0_io_TOP_AXI_ARVALID = io_TOP_AXI_ARVALID;
  assign mags_0_io_TOP_AXI_ARREADY = io_TOP_AXI_ARREADY;
  assign mags_0_io_TOP_AXI_WDATA = io_TOP_AXI_WDATA;
  assign mags_0_io_TOP_AXI_WSTRB = io_TOP_AXI_WSTRB;
  assign mags_0_io_TOP_AXI_WVALID = io_TOP_AXI_WVALID;
  assign mags_0_io_TOP_AXI_WREADY = io_TOP_AXI_WREADY;
  assign mags_0_io_TOP_AXI_RVALID = io_TOP_AXI_RVALID;
  assign mags_0_io_TOP_AXI_RREADY = io_TOP_AXI_RREADY;
  assign mags_0_io_TOP_AXI_BVALID = io_TOP_AXI_BVALID;
  assign mags_0_io_TOP_AXI_BREADY = io_TOP_AXI_BREADY;
  assign mags_0_io_DWIDTH_AXI_AWADDR = io_DWIDTH_AXI_AWADDR;
  assign mags_0_io_DWIDTH_AXI_AWLEN = io_DWIDTH_AXI_AWLEN;
  assign mags_0_io_DWIDTH_AXI_AWVALID = io_DWIDTH_AXI_AWVALID;
  assign mags_0_io_DWIDTH_AXI_AWREADY = io_DWIDTH_AXI_AWREADY;
  assign mags_0_io_DWIDTH_AXI_ARADDR = io_DWIDTH_AXI_ARADDR;
  assign mags_0_io_DWIDTH_AXI_ARLEN = io_DWIDTH_AXI_ARLEN;
  assign mags_0_io_DWIDTH_AXI_ARSIZE = io_DWIDTH_AXI_ARSIZE;
  assign mags_0_io_DWIDTH_AXI_ARBURST = io_DWIDTH_AXI_ARBURST;
  assign mags_0_io_DWIDTH_AXI_ARVALID = io_DWIDTH_AXI_ARVALID;
  assign mags_0_io_DWIDTH_AXI_ARREADY = io_DWIDTH_AXI_ARREADY;
  assign mags_0_io_DWIDTH_AXI_WDATA = io_DWIDTH_AXI_WDATA;
  assign mags_0_io_DWIDTH_AXI_WSTRB = io_DWIDTH_AXI_WSTRB;
  assign mags_0_io_DWIDTH_AXI_WVALID = io_DWIDTH_AXI_WVALID;
  assign mags_0_io_DWIDTH_AXI_WREADY = io_DWIDTH_AXI_WREADY;
  assign mags_0_io_DWIDTH_AXI_RVALID = io_DWIDTH_AXI_RVALID;
  assign mags_0_io_DWIDTH_AXI_RREADY = io_DWIDTH_AXI_RREADY;
  assign mags_0_io_DWIDTH_AXI_BVALID = io_DWIDTH_AXI_BVALID;
  assign mags_0_io_DWIDTH_AXI_BREADY = io_DWIDTH_AXI_BREADY;
  assign mags_0_clock = clock;
  assign mags_0_reset = localReset;
  assign mags_1_io_enable = localEnable;
  assign mags_1_io_reset = localReset;
  assign mags_1_io_app_loads_0_cmd_valid = io_memStreams_loads_2_cmd_valid;
  assign mags_1_io_app_loads_0_cmd_bits_addr = io_memStreams_loads_2_cmd_bits_addr;
  assign mags_1_io_app_loads_0_cmd_bits_isWr = io_memStreams_loads_2_cmd_bits_isWr;
  assign mags_1_io_app_loads_0_cmd_bits_size = io_memStreams_loads_2_cmd_bits_size;
  assign mags_1_io_app_loads_0_rdata_ready = io_memStreams_loads_2_rdata_ready;
  assign mags_1_io_dram_cmd_ready = io_dram_1_cmd_ready;
  assign mags_1_io_dram_wdata_ready = io_dram_1_wdata_ready;
  assign mags_1_io_dram_rresp_valid = io_dram_1_rresp_valid;
  assign mags_1_io_dram_rresp_bits_rdata_0 = io_dram_1_rresp_bits_rdata_0;
  assign mags_1_io_dram_rresp_bits_rdata_1 = io_dram_1_rresp_bits_rdata_1;
  assign mags_1_io_dram_rresp_bits_rdata_2 = io_dram_1_rresp_bits_rdata_2;
  assign mags_1_io_dram_rresp_bits_rdata_3 = io_dram_1_rresp_bits_rdata_3;
  assign mags_1_io_dram_rresp_bits_rdata_4 = io_dram_1_rresp_bits_rdata_4;
  assign mags_1_io_dram_rresp_bits_rdata_5 = io_dram_1_rresp_bits_rdata_5;
  assign mags_1_io_dram_rresp_bits_rdata_6 = io_dram_1_rresp_bits_rdata_6;
  assign mags_1_io_dram_rresp_bits_rdata_7 = io_dram_1_rresp_bits_rdata_7;
  assign mags_1_io_dram_rresp_bits_rdata_8 = io_dram_1_rresp_bits_rdata_8;
  assign mags_1_io_dram_rresp_bits_rdata_9 = io_dram_1_rresp_bits_rdata_9;
  assign mags_1_io_dram_rresp_bits_rdata_10 = io_dram_1_rresp_bits_rdata_10;
  assign mags_1_io_dram_rresp_bits_rdata_11 = io_dram_1_rresp_bits_rdata_11;
  assign mags_1_io_dram_rresp_bits_rdata_12 = io_dram_1_rresp_bits_rdata_12;
  assign mags_1_io_dram_rresp_bits_rdata_13 = io_dram_1_rresp_bits_rdata_13;
  assign mags_1_io_dram_rresp_bits_rdata_14 = io_dram_1_rresp_bits_rdata_14;
  assign mags_1_io_dram_rresp_bits_rdata_15 = io_dram_1_rresp_bits_rdata_15;
  assign mags_1_io_dram_rresp_bits_tag_streamId = io_dram_1_rresp_bits_tag_streamId;
  assign mags_1_io_dram_wresp_valid = io_dram_1_wresp_valid;
  assign mags_1_io_dram_wresp_bits_tag_streamId = io_dram_1_wresp_bits_tag_streamId;
  assign mags_1_clock = clock;
  assign mags_1_reset = localReset;
  assign mags_2_io_enable = localEnable;
  assign mags_2_io_reset = localReset;
  assign mags_2_io_app_loads_0_cmd_valid = io_memStreams_loads_1_cmd_valid;
  assign mags_2_io_app_loads_0_cmd_bits_addr = io_memStreams_loads_1_cmd_bits_addr;
  assign mags_2_io_app_loads_0_cmd_bits_isWr = io_memStreams_loads_1_cmd_bits_isWr;
  assign mags_2_io_app_loads_0_cmd_bits_size = io_memStreams_loads_1_cmd_bits_size;
  assign mags_2_io_app_loads_0_rdata_ready = io_memStreams_loads_1_rdata_ready;
  assign mags_2_io_dram_cmd_ready = io_dram_2_cmd_ready;
  assign mags_2_io_dram_wdata_ready = io_dram_2_wdata_ready;
  assign mags_2_io_dram_rresp_valid = io_dram_2_rresp_valid;
  assign mags_2_io_dram_rresp_bits_rdata_0 = io_dram_2_rresp_bits_rdata_0;
  assign mags_2_io_dram_rresp_bits_rdata_1 = io_dram_2_rresp_bits_rdata_1;
  assign mags_2_io_dram_rresp_bits_rdata_2 = io_dram_2_rresp_bits_rdata_2;
  assign mags_2_io_dram_rresp_bits_rdata_3 = io_dram_2_rresp_bits_rdata_3;
  assign mags_2_io_dram_rresp_bits_rdata_4 = io_dram_2_rresp_bits_rdata_4;
  assign mags_2_io_dram_rresp_bits_rdata_5 = io_dram_2_rresp_bits_rdata_5;
  assign mags_2_io_dram_rresp_bits_rdata_6 = io_dram_2_rresp_bits_rdata_6;
  assign mags_2_io_dram_rresp_bits_rdata_7 = io_dram_2_rresp_bits_rdata_7;
  assign mags_2_io_dram_rresp_bits_rdata_8 = io_dram_2_rresp_bits_rdata_8;
  assign mags_2_io_dram_rresp_bits_rdata_9 = io_dram_2_rresp_bits_rdata_9;
  assign mags_2_io_dram_rresp_bits_rdata_10 = io_dram_2_rresp_bits_rdata_10;
  assign mags_2_io_dram_rresp_bits_rdata_11 = io_dram_2_rresp_bits_rdata_11;
  assign mags_2_io_dram_rresp_bits_rdata_12 = io_dram_2_rresp_bits_rdata_12;
  assign mags_2_io_dram_rresp_bits_rdata_13 = io_dram_2_rresp_bits_rdata_13;
  assign mags_2_io_dram_rresp_bits_rdata_14 = io_dram_2_rresp_bits_rdata_14;
  assign mags_2_io_dram_rresp_bits_rdata_15 = io_dram_2_rresp_bits_rdata_15;
  assign mags_2_io_dram_rresp_bits_tag_streamId = io_dram_2_rresp_bits_tag_streamId;
  assign mags_2_io_dram_wresp_valid = io_dram_2_wresp_valid;
  assign mags_2_io_dram_wresp_bits_tag_streamId = io_dram_2_wresp_bits_tag_streamId;
  assign mags_2_clock = clock;
  assign mags_2_reset = localReset;
  assign mags_3_io_enable = localEnable;
  assign mags_3_io_reset = localReset;
  assign mags_3_io_app_loads_0_cmd_valid = io_memStreams_loads_0_cmd_valid;
  assign mags_3_io_app_loads_0_cmd_bits_addr = io_memStreams_loads_0_cmd_bits_addr;
  assign mags_3_io_app_loads_0_cmd_bits_isWr = io_memStreams_loads_0_cmd_bits_isWr;
  assign mags_3_io_app_loads_0_cmd_bits_size = io_memStreams_loads_0_cmd_bits_size;
  assign mags_3_io_app_loads_0_rdata_ready = io_memStreams_loads_0_rdata_ready;
  assign mags_3_io_dram_cmd_ready = io_dram_3_cmd_ready;
  assign mags_3_io_dram_wdata_ready = io_dram_3_wdata_ready;
  assign mags_3_io_dram_rresp_valid = io_dram_3_rresp_valid;
  assign mags_3_io_dram_rresp_bits_rdata_0 = io_dram_3_rresp_bits_rdata_0;
  assign mags_3_io_dram_rresp_bits_rdata_1 = io_dram_3_rresp_bits_rdata_1;
  assign mags_3_io_dram_rresp_bits_rdata_2 = io_dram_3_rresp_bits_rdata_2;
  assign mags_3_io_dram_rresp_bits_rdata_3 = io_dram_3_rresp_bits_rdata_3;
  assign mags_3_io_dram_rresp_bits_rdata_4 = io_dram_3_rresp_bits_rdata_4;
  assign mags_3_io_dram_rresp_bits_rdata_5 = io_dram_3_rresp_bits_rdata_5;
  assign mags_3_io_dram_rresp_bits_rdata_6 = io_dram_3_rresp_bits_rdata_6;
  assign mags_3_io_dram_rresp_bits_rdata_7 = io_dram_3_rresp_bits_rdata_7;
  assign mags_3_io_dram_rresp_bits_rdata_8 = io_dram_3_rresp_bits_rdata_8;
  assign mags_3_io_dram_rresp_bits_rdata_9 = io_dram_3_rresp_bits_rdata_9;
  assign mags_3_io_dram_rresp_bits_rdata_10 = io_dram_3_rresp_bits_rdata_10;
  assign mags_3_io_dram_rresp_bits_rdata_11 = io_dram_3_rresp_bits_rdata_11;
  assign mags_3_io_dram_rresp_bits_rdata_12 = io_dram_3_rresp_bits_rdata_12;
  assign mags_3_io_dram_rresp_bits_rdata_13 = io_dram_3_rresp_bits_rdata_13;
  assign mags_3_io_dram_rresp_bits_rdata_14 = io_dram_3_rresp_bits_rdata_14;
  assign mags_3_io_dram_rresp_bits_rdata_15 = io_dram_3_rresp_bits_rdata_15;
  assign mags_3_io_dram_rresp_bits_tag_streamId = io_dram_3_rresp_bits_tag_streamId;
  assign mags_3_io_dram_wresp_valid = io_dram_3_wresp_valid;
  assign mags_3_io_dram_wresp_bits_tag_streamId = io_dram_3_wresp_bits_tag_streamId;
  assign mags_3_clock = clock;
  assign mags_3_reset = localReset;
  assign regs_io_raddr = io_raddr;
  assign regs_io_wen = io_wen;
  assign regs_io_waddr = io_waddr;
  assign regs_io_wdata = io_wdata;
  assign regs_io_reset = localReset;
  assign regs_io_argOuts_0_valid = status_valid;
  assign regs_io_argOuts_0_bits = status_bits;
  assign regs_io_argOuts_1_valid = io_argOuts_0_valid;
  assign regs_io_argOuts_1_bits = io_argOuts_0_bits;
  assign regs_io_argOuts_2_bits = {{32'd0}, mags_0_io_debugSignals_0};
  assign regs_io_argOuts_3_bits = {{32'd0}, mags_0_io_debugSignals_1};
  assign regs_io_argOuts_4_bits = {{32'd0}, mags_0_io_debugSignals_2};
  assign regs_io_argOuts_5_bits = {{32'd0}, mags_0_io_debugSignals_3};
  assign regs_io_argOuts_6_bits = {{32'd0}, mags_0_io_debugSignals_4};
  assign regs_io_argOuts_7_bits = {{32'd0}, mags_0_io_debugSignals_5};
  assign regs_io_argOuts_8_bits = {{32'd0}, mags_0_io_debugSignals_6};
  assign regs_io_argOuts_9_bits = {{32'd0}, mags_0_io_debugSignals_7};
  assign regs_io_argOuts_10_bits = {{32'd0}, mags_0_io_debugSignals_8};
  assign regs_io_argOuts_11_bits = {{32'd0}, mags_0_io_debugSignals_9};
  assign regs_io_argOuts_12_bits = {{32'd0}, mags_0_io_debugSignals_10};
  assign regs_io_argOuts_13_bits = {{32'd0}, mags_0_io_debugSignals_11};
  assign regs_io_argOuts_14_bits = {{32'd0}, mags_0_io_debugSignals_12};
  assign regs_io_argOuts_15_bits = {{32'd0}, mags_0_io_debugSignals_13};
  assign regs_io_argOuts_16_bits = {{32'd0}, mags_0_io_debugSignals_14};
  assign regs_io_argOuts_17_bits = {{32'd0}, mags_0_io_debugSignals_15};
  assign regs_io_argOuts_18_bits = {{32'd0}, mags_0_io_debugSignals_16};
  assign regs_io_argOuts_19_bits = {{32'd0}, mags_0_io_debugSignals_17};
  assign regs_io_argOuts_20_bits = {{32'd0}, mags_0_io_debugSignals_18};
  assign regs_io_argOuts_21_bits = {{32'd0}, mags_0_io_debugSignals_19};
  assign regs_io_argOuts_22_bits = {{32'd0}, mags_0_io_debugSignals_20};
  assign regs_io_argOuts_23_bits = {{32'd0}, mags_0_io_debugSignals_21};
  assign regs_io_argOuts_24_bits = {{32'd0}, mags_0_io_debugSignals_22};
  assign regs_io_argOuts_25_bits = {{32'd0}, mags_0_io_debugSignals_23};
  assign regs_io_argOuts_26_bits = {{32'd0}, mags_0_io_debugSignals_24};
  assign regs_io_argOuts_27_bits = {{32'd0}, mags_0_io_debugSignals_25};
  assign regs_io_argOuts_28_bits = {{32'd0}, mags_0_io_debugSignals_26};
  assign regs_io_argOuts_29_bits = {{32'd0}, mags_0_io_debugSignals_27};
  assign regs_io_argOuts_30_bits = {{32'd0}, mags_0_io_debugSignals_28};
  assign regs_io_argOuts_31_bits = {{32'd0}, mags_0_io_debugSignals_29};
  assign regs_io_argOuts_32_bits = {{32'd0}, mags_0_io_debugSignals_30};
  assign regs_io_argOuts_33_bits = {{32'd0}, mags_0_io_debugSignals_31};
  assign regs_io_argOuts_34_bits = {{32'd0}, mags_0_io_debugSignals_32};
  assign regs_io_argOuts_35_bits = {{32'd0}, mags_0_io_debugSignals_33};
  assign regs_io_argOuts_36_bits = {{32'd0}, mags_0_io_debugSignals_34};
  assign regs_io_argOuts_37_bits = {{32'd0}, mags_0_io_debugSignals_35};
  assign regs_io_argOuts_38_bits = {{32'd0}, mags_0_io_debugSignals_36};
  assign regs_io_argOuts_39_bits = {{32'd0}, mags_0_io_debugSignals_37};
  assign regs_io_argOuts_40_bits = {{32'd0}, mags_0_io_debugSignals_38};
  assign regs_io_argOuts_41_bits = {{32'd0}, mags_0_io_debugSignals_39};
  assign regs_io_argOuts_42_bits = {{32'd0}, mags_0_io_debugSignals_40};
  assign regs_io_argOuts_43_bits = {{32'd0}, mags_0_io_debugSignals_41};
  assign regs_io_argOuts_44_bits = {{32'd0}, mags_0_io_debugSignals_42};
  assign regs_io_argOuts_45_bits = {{32'd0}, mags_0_io_debugSignals_43};
  assign regs_io_argOuts_46_bits = {{32'd0}, mags_0_io_debugSignals_44};
  assign regs_io_argOuts_47_bits = {{32'd0}, mags_0_io_debugSignals_45};
  assign regs_io_argOuts_48_bits = {{32'd0}, mags_0_io_debugSignals_46};
  assign regs_io_argOuts_49_bits = {{32'd0}, mags_0_io_debugSignals_47};
  assign regs_io_argOuts_50_bits = {{32'd0}, mags_0_io_debugSignals_48};
  assign regs_io_argOuts_51_bits = {{32'd0}, mags_0_io_debugSignals_49};
  assign regs_io_argOuts_52_bits = {{32'd0}, mags_0_io_debugSignals_50};
  assign regs_io_argOuts_53_bits = {{32'd0}, mags_0_io_debugSignals_51};
  assign regs_io_argOuts_54_bits = {{32'd0}, mags_0_io_debugSignals_52};
  assign regs_io_argOuts_55_bits = {{32'd0}, mags_0_io_debugSignals_53};
  assign regs_io_argOuts_56_bits = {{32'd0}, mags_0_io_debugSignals_54};
  assign regs_io_argOuts_57_bits = {{32'd0}, mags_0_io_debugSignals_55};
  assign regs_io_argOuts_58_bits = {{32'd0}, mags_0_io_debugSignals_56};
  assign regs_io_argOuts_59_bits = {{32'd0}, mags_0_io_debugSignals_57};
  assign regs_io_argOuts_60_bits = {{32'd0}, mags_0_io_debugSignals_58};
  assign regs_io_argOuts_61_bits = {{32'd0}, mags_0_io_debugSignals_59};
  assign regs_io_argOuts_62_bits = {{32'd0}, mags_0_io_debugSignals_60};
  assign regs_io_argOuts_63_bits = {{32'd0}, mags_0_io_debugSignals_61};
  assign regs_io_argOuts_64_bits = {{32'd0}, mags_0_io_debugSignals_62};
  assign regs_io_argOuts_65_bits = {{32'd0}, mags_0_io_debugSignals_63};
  assign regs_io_argOuts_66_bits = {{32'd0}, mags_0_io_debugSignals_64};
  assign regs_io_argOuts_67_bits = {{32'd0}, mags_0_io_debugSignals_65};
  assign regs_io_argOuts_68_bits = {{32'd0}, mags_0_io_debugSignals_66};
  assign regs_io_argOuts_69_bits = {{32'd0}, mags_0_io_debugSignals_67};
  assign regs_io_argOuts_70_bits = {{32'd0}, mags_0_io_debugSignals_68};
  assign regs_io_argOuts_71_bits = {{32'd0}, mags_0_io_debugSignals_69};
  assign regs_io_argOuts_72_bits = {{32'd0}, mags_0_io_debugSignals_70};
  assign regs_io_argOuts_73_bits = {{32'd0}, mags_0_io_debugSignals_71};
  assign regs_io_argOuts_74_bits = {{32'd0}, mags_0_io_debugSignals_72};
  assign regs_io_argOuts_75_bits = {{32'd0}, mags_0_io_debugSignals_73};
  assign regs_io_argOuts_76_bits = {{32'd0}, mags_0_io_debugSignals_74};
  assign regs_io_argOuts_77_bits = {{32'd0}, mags_0_io_debugSignals_75};
  assign regs_io_argOuts_78_bits = {{32'd0}, mags_0_io_debugSignals_76};
  assign regs_io_argOuts_79_bits = {{32'd0}, mags_0_io_debugSignals_77};
  assign regs_io_argOuts_80_bits = {{32'd0}, mags_0_io_debugSignals_78};
  assign regs_io_argOuts_81_bits = {{32'd0}, mags_0_io_debugSignals_79};
  assign regs_io_argOuts_82_bits = {{32'd0}, mags_0_io_debugSignals_80};
  assign regs_io_argOuts_83_bits = {{32'd0}, mags_0_io_debugSignals_81};
  assign regs_io_argOuts_84_bits = {{32'd0}, mags_0_io_debugSignals_82};
  assign regs_io_argOuts_85_bits = {{32'd0}, mags_0_io_debugSignals_83};
  assign regs_io_argOuts_86_bits = {{32'd0}, mags_0_io_debugSignals_84};
  assign regs_io_argOuts_87_bits = {{32'd0}, mags_0_io_debugSignals_85};
  assign regs_io_argOuts_88_bits = {{32'd0}, mags_0_io_debugSignals_86};
  assign regs_io_argOuts_89_bits = {{32'd0}, mags_0_io_debugSignals_87};
  assign regs_io_argOuts_90_bits = {{32'd0}, mags_0_io_debugSignals_88};
  assign regs_io_argOuts_91_bits = {{32'd0}, mags_0_io_debugSignals_89};
  assign regs_io_argOuts_92_bits = {{32'd0}, mags_0_io_debugSignals_90};
  assign regs_io_argOuts_93_bits = {{32'd0}, mags_0_io_debugSignals_91};
  assign regs_io_argOuts_94_bits = {{32'd0}, mags_0_io_debugSignals_92};
  assign regs_io_argOuts_95_bits = {{32'd0}, mags_0_io_debugSignals_93};
  assign regs_io_argOuts_96_bits = {{32'd0}, mags_0_io_debugSignals_94};
  assign regs_io_argOuts_97_bits = {{32'd0}, mags_0_io_debugSignals_95};
  assign regs_io_argOuts_98_bits = {{32'd0}, mags_0_io_debugSignals_96};
  assign regs_io_argOuts_99_bits = {{32'd0}, mags_0_io_debugSignals_97};
  assign regs_io_argOuts_100_bits = {{32'd0}, mags_0_io_debugSignals_98};
  assign regs_io_argOuts_101_bits = {{32'd0}, mags_0_io_debugSignals_99};
  assign regs_io_argOuts_102_bits = {{32'd0}, mags_0_io_debugSignals_100};
  assign regs_io_argOuts_103_bits = {{32'd0}, mags_0_io_debugSignals_101};
  assign regs_io_argOuts_104_bits = {{32'd0}, mags_0_io_debugSignals_102};
  assign regs_io_argOuts_105_bits = {{32'd0}, mags_0_io_debugSignals_103};
  assign regs_io_argOuts_106_bits = {{32'd0}, mags_0_io_debugSignals_104};
  assign regs_io_argOuts_107_bits = {{32'd0}, mags_0_io_debugSignals_105};
  assign regs_io_argOuts_108_bits = {{32'd0}, mags_0_io_debugSignals_106};
  assign regs_io_argOuts_109_bits = {{32'd0}, mags_0_io_debugSignals_107};
  assign regs_clock = clock;
  assign regs_reset = reset;
  assign timeoutCtr_io_enable = localEnable;
  assign timeoutCtr_clock = clock;
  assign timeoutCtr_reset = reset;
  assign depulser_io_in = _T_726;
  assign depulser_io_rst = _T_727[0];
  assign depulser_clock = clock;
  assign depulser_reset = reset;
  assign status_valid = depulser_io_out;
  assign status_bits = {{62'd0}, _T_740};
endmodule
module AXI4LiteToRFBridge(
  input         clock,
  input         reset,
  input  [31:0] io_S_AXI_AWADDR,
  input  [2:0]  io_S_AXI_AWPROT,
  input         io_S_AXI_AWVALID,
  output        io_S_AXI_AWREADY,
  input  [31:0] io_S_AXI_ARADDR,
  input  [2:0]  io_S_AXI_ARPROT,
  input         io_S_AXI_ARVALID,
  output        io_S_AXI_ARREADY,
  input  [31:0] io_S_AXI_WDATA,
  input  [3:0]  io_S_AXI_WSTRB,
  input         io_S_AXI_WVALID,
  output        io_S_AXI_WREADY,
  output [31:0] io_S_AXI_RDATA,
  output [1:0]  io_S_AXI_RRESP,
  output        io_S_AXI_RVALID,
  input         io_S_AXI_RREADY,
  output [1:0]  io_S_AXI_BRESP,
  output        io_S_AXI_BVALID,
  input         io_S_AXI_BREADY,
  output [31:0] io_raddr,
  output        io_wen,
  output [31:0] io_waddr,
  output [31:0] io_wdata,
  input  [31:0] io_rdata
);
  wire [31:0] d_rf_rdata;
  wire [31:0] d_rf_wdata;
  wire [31:0] d_rf_waddr;
  wire  d_rf_wen;
  wire [31:0] d_rf_raddr;
  wire  d_S_AXI_ARESETN;
  wire  d_S_AXI_ACLK;
  wire [31:0] d_S_AXI_AWADDR;
  wire [2:0] d_S_AXI_AWPROT;
  wire  d_S_AXI_AWVALID;
  wire  d_S_AXI_AWREADY;
  wire [31:0] d_S_AXI_ARADDR;
  wire [2:0] d_S_AXI_ARPROT;
  wire  d_S_AXI_ARVALID;
  wire  d_S_AXI_ARREADY;
  wire [31:0] d_S_AXI_WDATA;
  wire [3:0] d_S_AXI_WSTRB;
  wire  d_S_AXI_WVALID;
  wire  d_S_AXI_WREADY;
  wire [31:0] d_S_AXI_RDATA;
  wire [1:0] d_S_AXI_RRESP;
  wire  d_S_AXI_RVALID;
  wire  d_S_AXI_RREADY;
  wire [1:0] d_S_AXI_BRESP;
  wire  d_S_AXI_BVALID;
  wire  d_S_AXI_BREADY;
  wire  _T_47;
  AXI4LiteToRFBridgeVerilog d (
    .rf_rdata(d_rf_rdata),
    .rf_wdata(d_rf_wdata),
    .rf_waddr(d_rf_waddr),
    .rf_wen(d_rf_wen),
    .rf_raddr(d_rf_raddr),
    .S_AXI_ARESETN(d_S_AXI_ARESETN),
    .S_AXI_ACLK(d_S_AXI_ACLK),
    .S_AXI_AWADDR(d_S_AXI_AWADDR),
    .S_AXI_AWPROT(d_S_AXI_AWPROT),
    .S_AXI_AWVALID(d_S_AXI_AWVALID),
    .S_AXI_AWREADY(d_S_AXI_AWREADY),
    .S_AXI_ARADDR(d_S_AXI_ARADDR),
    .S_AXI_ARPROT(d_S_AXI_ARPROT),
    .S_AXI_ARVALID(d_S_AXI_ARVALID),
    .S_AXI_ARREADY(d_S_AXI_ARREADY),
    .S_AXI_WDATA(d_S_AXI_WDATA),
    .S_AXI_WSTRB(d_S_AXI_WSTRB),
    .S_AXI_WVALID(d_S_AXI_WVALID),
    .S_AXI_WREADY(d_S_AXI_WREADY),
    .S_AXI_RDATA(d_S_AXI_RDATA),
    .S_AXI_RRESP(d_S_AXI_RRESP),
    .S_AXI_RVALID(d_S_AXI_RVALID),
    .S_AXI_RREADY(d_S_AXI_RREADY),
    .S_AXI_BRESP(d_S_AXI_BRESP),
    .S_AXI_BVALID(d_S_AXI_BVALID),
    .S_AXI_BREADY(d_S_AXI_BREADY)
  );
  assign _T_47 = ~ reset;
  assign io_S_AXI_AWREADY = d_S_AXI_AWREADY;
  assign io_S_AXI_ARREADY = d_S_AXI_ARREADY;
  assign io_S_AXI_WREADY = d_S_AXI_WREADY;
  assign io_S_AXI_RDATA = d_S_AXI_RDATA;
  assign io_S_AXI_RRESP = d_S_AXI_RRESP;
  assign io_S_AXI_RVALID = d_S_AXI_RVALID;
  assign io_S_AXI_BRESP = d_S_AXI_BRESP;
  assign io_S_AXI_BVALID = d_S_AXI_BVALID;
  assign io_raddr = d_rf_raddr;
  assign io_wen = d_rf_wen;
  assign io_waddr = d_rf_waddr;
  assign io_wdata = d_rf_wdata;
  assign d_rf_rdata = io_rdata;
  assign d_S_AXI_ARESETN = _T_47;
  assign d_S_AXI_ACLK = clock;
  assign d_S_AXI_AWADDR = io_S_AXI_AWADDR;
  assign d_S_AXI_AWPROT = io_S_AXI_AWPROT;
  assign d_S_AXI_AWVALID = io_S_AXI_AWVALID;
  assign d_S_AXI_ARADDR = io_S_AXI_ARADDR;
  assign d_S_AXI_ARPROT = io_S_AXI_ARPROT;
  assign d_S_AXI_ARVALID = io_S_AXI_ARVALID;
  assign d_S_AXI_WDATA = io_S_AXI_WDATA;
  assign d_S_AXI_WSTRB = io_S_AXI_WSTRB;
  assign d_S_AXI_WVALID = io_S_AXI_WVALID;
  assign d_S_AXI_RREADY = io_S_AXI_RREADY;
  assign d_S_AXI_BREADY = io_S_AXI_BREADY;
endmodule
module MAGToAXI4Bridge(
  output         io_in_cmd_ready,
  input          io_in_cmd_valid,
  input  [63:0]  io_in_cmd_bits_addr,
  input  [31:0]  io_in_cmd_bits_size,
  input          io_in_cmd_bits_isWr,
  input  [25:0]  io_in_cmd_bits_tag_uid,
  input  [5:0]   io_in_cmd_bits_tag_streamId,
  output         io_in_wdata_ready,
  input          io_in_wdata_valid,
  input  [31:0]  io_in_wdata_bits_wdata_0,
  input  [31:0]  io_in_wdata_bits_wdata_1,
  input  [31:0]  io_in_wdata_bits_wdata_2,
  input  [31:0]  io_in_wdata_bits_wdata_3,
  input  [31:0]  io_in_wdata_bits_wdata_4,
  input  [31:0]  io_in_wdata_bits_wdata_5,
  input  [31:0]  io_in_wdata_bits_wdata_6,
  input  [31:0]  io_in_wdata_bits_wdata_7,
  input  [31:0]  io_in_wdata_bits_wdata_8,
  input  [31:0]  io_in_wdata_bits_wdata_9,
  input  [31:0]  io_in_wdata_bits_wdata_10,
  input  [31:0]  io_in_wdata_bits_wdata_11,
  input  [31:0]  io_in_wdata_bits_wdata_12,
  input  [31:0]  io_in_wdata_bits_wdata_13,
  input  [31:0]  io_in_wdata_bits_wdata_14,
  input  [31:0]  io_in_wdata_bits_wdata_15,
  input          io_in_wdata_bits_wstrb_0,
  input          io_in_wdata_bits_wstrb_1,
  input          io_in_wdata_bits_wstrb_2,
  input          io_in_wdata_bits_wstrb_3,
  input          io_in_wdata_bits_wstrb_4,
  input          io_in_wdata_bits_wstrb_5,
  input          io_in_wdata_bits_wstrb_6,
  input          io_in_wdata_bits_wstrb_7,
  input          io_in_wdata_bits_wstrb_8,
  input          io_in_wdata_bits_wstrb_9,
  input          io_in_wdata_bits_wstrb_10,
  input          io_in_wdata_bits_wstrb_11,
  input          io_in_wdata_bits_wstrb_12,
  input          io_in_wdata_bits_wstrb_13,
  input          io_in_wdata_bits_wstrb_14,
  input          io_in_wdata_bits_wstrb_15,
  input          io_in_wdata_bits_wstrb_16,
  input          io_in_wdata_bits_wstrb_17,
  input          io_in_wdata_bits_wstrb_18,
  input          io_in_wdata_bits_wstrb_19,
  input          io_in_wdata_bits_wstrb_20,
  input          io_in_wdata_bits_wstrb_21,
  input          io_in_wdata_bits_wstrb_22,
  input          io_in_wdata_bits_wstrb_23,
  input          io_in_wdata_bits_wstrb_24,
  input          io_in_wdata_bits_wstrb_25,
  input          io_in_wdata_bits_wstrb_26,
  input          io_in_wdata_bits_wstrb_27,
  input          io_in_wdata_bits_wstrb_28,
  input          io_in_wdata_bits_wstrb_29,
  input          io_in_wdata_bits_wstrb_30,
  input          io_in_wdata_bits_wstrb_31,
  input          io_in_wdata_bits_wstrb_32,
  input          io_in_wdata_bits_wstrb_33,
  input          io_in_wdata_bits_wstrb_34,
  input          io_in_wdata_bits_wstrb_35,
  input          io_in_wdata_bits_wstrb_36,
  input          io_in_wdata_bits_wstrb_37,
  input          io_in_wdata_bits_wstrb_38,
  input          io_in_wdata_bits_wstrb_39,
  input          io_in_wdata_bits_wstrb_40,
  input          io_in_wdata_bits_wstrb_41,
  input          io_in_wdata_bits_wstrb_42,
  input          io_in_wdata_bits_wstrb_43,
  input          io_in_wdata_bits_wstrb_44,
  input          io_in_wdata_bits_wstrb_45,
  input          io_in_wdata_bits_wstrb_46,
  input          io_in_wdata_bits_wstrb_47,
  input          io_in_wdata_bits_wstrb_48,
  input          io_in_wdata_bits_wstrb_49,
  input          io_in_wdata_bits_wstrb_50,
  input          io_in_wdata_bits_wstrb_51,
  input          io_in_wdata_bits_wstrb_52,
  input          io_in_wdata_bits_wstrb_53,
  input          io_in_wdata_bits_wstrb_54,
  input          io_in_wdata_bits_wstrb_55,
  input          io_in_wdata_bits_wstrb_56,
  input          io_in_wdata_bits_wstrb_57,
  input          io_in_wdata_bits_wstrb_58,
  input          io_in_wdata_bits_wstrb_59,
  input          io_in_wdata_bits_wstrb_60,
  input          io_in_wdata_bits_wstrb_61,
  input          io_in_wdata_bits_wstrb_62,
  input          io_in_wdata_bits_wstrb_63,
  input          io_in_rresp_ready,
  output         io_in_rresp_valid,
  output [31:0]  io_in_rresp_bits_rdata_0,
  output [31:0]  io_in_rresp_bits_rdata_1,
  output [31:0]  io_in_rresp_bits_rdata_2,
  output [31:0]  io_in_rresp_bits_rdata_3,
  output [31:0]  io_in_rresp_bits_rdata_4,
  output [31:0]  io_in_rresp_bits_rdata_5,
  output [31:0]  io_in_rresp_bits_rdata_6,
  output [31:0]  io_in_rresp_bits_rdata_7,
  output [31:0]  io_in_rresp_bits_rdata_8,
  output [31:0]  io_in_rresp_bits_rdata_9,
  output [31:0]  io_in_rresp_bits_rdata_10,
  output [31:0]  io_in_rresp_bits_rdata_11,
  output [31:0]  io_in_rresp_bits_rdata_12,
  output [31:0]  io_in_rresp_bits_rdata_13,
  output [31:0]  io_in_rresp_bits_rdata_14,
  output [31:0]  io_in_rresp_bits_rdata_15,
  output [5:0]   io_in_rresp_bits_tag_streamId,
  input          io_in_wresp_ready,
  output         io_in_wresp_valid,
  output [5:0]   io_in_wresp_bits_tag_streamId,
  output [31:0]  io_M_AXI_AWID,
  output [31:0]  io_M_AXI_AWADDR,
  output [7:0]   io_M_AXI_AWLEN,
  output         io_M_AXI_AWVALID,
  input          io_M_AXI_AWREADY,
  output [31:0]  io_M_AXI_ARID,
  output [31:0]  io_M_AXI_ARADDR,
  output [7:0]   io_M_AXI_ARLEN,
  output         io_M_AXI_ARVALID,
  input          io_M_AXI_ARREADY,
  output [511:0] io_M_AXI_WDATA,
  output [63:0]  io_M_AXI_WSTRB,
  output         io_M_AXI_WVALID,
  input          io_M_AXI_WREADY,
  input  [31:0]  io_M_AXI_RID,
  input  [511:0] io_M_AXI_RDATA,
  input          io_M_AXI_RVALID,
  output         io_M_AXI_RREADY,
  input  [31:0]  io_M_AXI_BID,
  input          io_M_AXI_BVALID,
  output         io_M_AXI_BREADY
);
  wire [31:0] id;
  wire [32:0] _T_137;
  wire [32:0] _T_138;
  wire [31:0] _T_139;
  wire  _T_146;
  wire  _T_147;
  wire  _T_148;
  wire  _T_159;
  wire [63:0] _T_160;
  wire [95:0] _T_161;
  wire [127:0] _T_162;
  wire [159:0] _T_163;
  wire [191:0] _T_164;
  wire [223:0] _T_165;
  wire [255:0] _T_166;
  wire [287:0] _T_167;
  wire [319:0] _T_168;
  wire [351:0] _T_169;
  wire [383:0] _T_170;
  wire [415:0] _T_171;
  wire [447:0] _T_172;
  wire [479:0] _T_173;
  wire [511:0] _T_174;
  wire [1:0] _T_175;
  wire [2:0] _T_176;
  wire [3:0] _T_177;
  wire [4:0] _T_178;
  wire [5:0] _T_179;
  wire [6:0] _T_180;
  wire [7:0] _T_181;
  wire [8:0] _T_182;
  wire [9:0] _T_183;
  wire [10:0] _T_184;
  wire [11:0] _T_185;
  wire [12:0] _T_186;
  wire [13:0] _T_187;
  wire [14:0] _T_188;
  wire [15:0] _T_189;
  wire [16:0] _T_190;
  wire [17:0] _T_191;
  wire [18:0] _T_192;
  wire [19:0] _T_193;
  wire [20:0] _T_194;
  wire [21:0] _T_195;
  wire [22:0] _T_196;
  wire [23:0] _T_197;
  wire [24:0] _T_198;
  wire [25:0] _T_199;
  wire [26:0] _T_200;
  wire [27:0] _T_201;
  wire [28:0] _T_202;
  wire [29:0] _T_203;
  wire [30:0] _T_204;
  wire [31:0] _T_205;
  wire [32:0] _T_206;
  wire [33:0] _T_207;
  wire [34:0] _T_208;
  wire [35:0] _T_209;
  wire [36:0] _T_210;
  wire [37:0] _T_211;
  wire [38:0] _T_212;
  wire [39:0] _T_213;
  wire [40:0] _T_214;
  wire [41:0] _T_215;
  wire [42:0] _T_216;
  wire [43:0] _T_217;
  wire [44:0] _T_218;
  wire [45:0] _T_219;
  wire [46:0] _T_220;
  wire [47:0] _T_221;
  wire [48:0] _T_222;
  wire [49:0] _T_223;
  wire [50:0] _T_224;
  wire [51:0] _T_225;
  wire [52:0] _T_226;
  wire [53:0] _T_227;
  wire [54:0] _T_228;
  wire [55:0] _T_229;
  wire [56:0] _T_230;
  wire [57:0] _T_231;
  wire [58:0] _T_232;
  wire [59:0] _T_233;
  wire [60:0] _T_234;
  wire [61:0] _T_235;
  wire [62:0] _T_236;
  wire [63:0] _T_237;
  wire [31:0] _T_238;
  wire [31:0] _T_239;
  wire [31:0] _T_240;
  wire [31:0] _T_241;
  wire [31:0] _T_242;
  wire [31:0] _T_243;
  wire [31:0] _T_244;
  wire [31:0] _T_245;
  wire [31:0] _T_246;
  wire [31:0] _T_247;
  wire [31:0] _T_248;
  wire [31:0] _T_249;
  wire [31:0] _T_250;
  wire [31:0] _T_251;
  wire [31:0] _T_252;
  wire [31:0] _T_253;
  wire [31:0] rdataAsVec_0;
  wire [31:0] rdataAsVec_1;
  wire [31:0] rdataAsVec_2;
  wire [31:0] rdataAsVec_3;
  wire [31:0] rdataAsVec_4;
  wire [31:0] rdataAsVec_5;
  wire [31:0] rdataAsVec_6;
  wire [31:0] rdataAsVec_7;
  wire [31:0] rdataAsVec_8;
  wire [31:0] rdataAsVec_9;
  wire [31:0] rdataAsVec_10;
  wire [31:0] rdataAsVec_11;
  wire [31:0] rdataAsVec_12;
  wire [31:0] rdataAsVec_13;
  wire [31:0] rdataAsVec_14;
  wire [31:0] rdataAsVec_15;
  wire [5:0] _T_276_streamId;
  wire [31:0] _T_278;
  wire [5:0] _T_279;
  wire [5:0] _T_283_streamId;
  wire [31:0] _T_285;
  wire [5:0] _T_286;
  assign id = {io_in_cmd_bits_tag_uid,io_in_cmd_bits_tag_streamId};
  assign _T_137 = io_in_cmd_bits_size - 32'h1;
  assign _T_138 = $unsigned(_T_137);
  assign _T_139 = _T_138[31:0];
  assign _T_146 = ~ io_in_cmd_bits_isWr;
  assign _T_147 = io_in_cmd_valid & _T_146;
  assign _T_148 = io_in_cmd_bits_isWr ? io_M_AXI_AWREADY : io_M_AXI_ARREADY;
  assign _T_159 = io_in_cmd_valid & io_in_cmd_bits_isWr;
  assign _T_160 = {io_in_wdata_bits_wdata_15,io_in_wdata_bits_wdata_14};
  assign _T_161 = {_T_160,io_in_wdata_bits_wdata_13};
  assign _T_162 = {_T_161,io_in_wdata_bits_wdata_12};
  assign _T_163 = {_T_162,io_in_wdata_bits_wdata_11};
  assign _T_164 = {_T_163,io_in_wdata_bits_wdata_10};
  assign _T_165 = {_T_164,io_in_wdata_bits_wdata_9};
  assign _T_166 = {_T_165,io_in_wdata_bits_wdata_8};
  assign _T_167 = {_T_166,io_in_wdata_bits_wdata_7};
  assign _T_168 = {_T_167,io_in_wdata_bits_wdata_6};
  assign _T_169 = {_T_168,io_in_wdata_bits_wdata_5};
  assign _T_170 = {_T_169,io_in_wdata_bits_wdata_4};
  assign _T_171 = {_T_170,io_in_wdata_bits_wdata_3};
  assign _T_172 = {_T_171,io_in_wdata_bits_wdata_2};
  assign _T_173 = {_T_172,io_in_wdata_bits_wdata_1};
  assign _T_174 = {_T_173,io_in_wdata_bits_wdata_0};
  assign _T_175 = {io_in_wdata_bits_wstrb_63,io_in_wdata_bits_wstrb_62};
  assign _T_176 = {_T_175,io_in_wdata_bits_wstrb_61};
  assign _T_177 = {_T_176,io_in_wdata_bits_wstrb_60};
  assign _T_178 = {_T_177,io_in_wdata_bits_wstrb_59};
  assign _T_179 = {_T_178,io_in_wdata_bits_wstrb_58};
  assign _T_180 = {_T_179,io_in_wdata_bits_wstrb_57};
  assign _T_181 = {_T_180,io_in_wdata_bits_wstrb_56};
  assign _T_182 = {_T_181,io_in_wdata_bits_wstrb_55};
  assign _T_183 = {_T_182,io_in_wdata_bits_wstrb_54};
  assign _T_184 = {_T_183,io_in_wdata_bits_wstrb_53};
  assign _T_185 = {_T_184,io_in_wdata_bits_wstrb_52};
  assign _T_186 = {_T_185,io_in_wdata_bits_wstrb_51};
  assign _T_187 = {_T_186,io_in_wdata_bits_wstrb_50};
  assign _T_188 = {_T_187,io_in_wdata_bits_wstrb_49};
  assign _T_189 = {_T_188,io_in_wdata_bits_wstrb_48};
  assign _T_190 = {_T_189,io_in_wdata_bits_wstrb_47};
  assign _T_191 = {_T_190,io_in_wdata_bits_wstrb_46};
  assign _T_192 = {_T_191,io_in_wdata_bits_wstrb_45};
  assign _T_193 = {_T_192,io_in_wdata_bits_wstrb_44};
  assign _T_194 = {_T_193,io_in_wdata_bits_wstrb_43};
  assign _T_195 = {_T_194,io_in_wdata_bits_wstrb_42};
  assign _T_196 = {_T_195,io_in_wdata_bits_wstrb_41};
  assign _T_197 = {_T_196,io_in_wdata_bits_wstrb_40};
  assign _T_198 = {_T_197,io_in_wdata_bits_wstrb_39};
  assign _T_199 = {_T_198,io_in_wdata_bits_wstrb_38};
  assign _T_200 = {_T_199,io_in_wdata_bits_wstrb_37};
  assign _T_201 = {_T_200,io_in_wdata_bits_wstrb_36};
  assign _T_202 = {_T_201,io_in_wdata_bits_wstrb_35};
  assign _T_203 = {_T_202,io_in_wdata_bits_wstrb_34};
  assign _T_204 = {_T_203,io_in_wdata_bits_wstrb_33};
  assign _T_205 = {_T_204,io_in_wdata_bits_wstrb_32};
  assign _T_206 = {_T_205,io_in_wdata_bits_wstrb_31};
  assign _T_207 = {_T_206,io_in_wdata_bits_wstrb_30};
  assign _T_208 = {_T_207,io_in_wdata_bits_wstrb_29};
  assign _T_209 = {_T_208,io_in_wdata_bits_wstrb_28};
  assign _T_210 = {_T_209,io_in_wdata_bits_wstrb_27};
  assign _T_211 = {_T_210,io_in_wdata_bits_wstrb_26};
  assign _T_212 = {_T_211,io_in_wdata_bits_wstrb_25};
  assign _T_213 = {_T_212,io_in_wdata_bits_wstrb_24};
  assign _T_214 = {_T_213,io_in_wdata_bits_wstrb_23};
  assign _T_215 = {_T_214,io_in_wdata_bits_wstrb_22};
  assign _T_216 = {_T_215,io_in_wdata_bits_wstrb_21};
  assign _T_217 = {_T_216,io_in_wdata_bits_wstrb_20};
  assign _T_218 = {_T_217,io_in_wdata_bits_wstrb_19};
  assign _T_219 = {_T_218,io_in_wdata_bits_wstrb_18};
  assign _T_220 = {_T_219,io_in_wdata_bits_wstrb_17};
  assign _T_221 = {_T_220,io_in_wdata_bits_wstrb_16};
  assign _T_222 = {_T_221,io_in_wdata_bits_wstrb_15};
  assign _T_223 = {_T_222,io_in_wdata_bits_wstrb_14};
  assign _T_224 = {_T_223,io_in_wdata_bits_wstrb_13};
  assign _T_225 = {_T_224,io_in_wdata_bits_wstrb_12};
  assign _T_226 = {_T_225,io_in_wdata_bits_wstrb_11};
  assign _T_227 = {_T_226,io_in_wdata_bits_wstrb_10};
  assign _T_228 = {_T_227,io_in_wdata_bits_wstrb_9};
  assign _T_229 = {_T_228,io_in_wdata_bits_wstrb_8};
  assign _T_230 = {_T_229,io_in_wdata_bits_wstrb_7};
  assign _T_231 = {_T_230,io_in_wdata_bits_wstrb_6};
  assign _T_232 = {_T_231,io_in_wdata_bits_wstrb_5};
  assign _T_233 = {_T_232,io_in_wdata_bits_wstrb_4};
  assign _T_234 = {_T_233,io_in_wdata_bits_wstrb_3};
  assign _T_235 = {_T_234,io_in_wdata_bits_wstrb_2};
  assign _T_236 = {_T_235,io_in_wdata_bits_wstrb_1};
  assign _T_237 = {_T_236,io_in_wdata_bits_wstrb_0};
  assign _T_238 = io_M_AXI_RDATA[511:480];
  assign _T_239 = io_M_AXI_RDATA[479:448];
  assign _T_240 = io_M_AXI_RDATA[447:416];
  assign _T_241 = io_M_AXI_RDATA[415:384];
  assign _T_242 = io_M_AXI_RDATA[383:352];
  assign _T_243 = io_M_AXI_RDATA[351:320];
  assign _T_244 = io_M_AXI_RDATA[319:288];
  assign _T_245 = io_M_AXI_RDATA[287:256];
  assign _T_246 = io_M_AXI_RDATA[255:224];
  assign _T_247 = io_M_AXI_RDATA[223:192];
  assign _T_248 = io_M_AXI_RDATA[191:160];
  assign _T_249 = io_M_AXI_RDATA[159:128];
  assign _T_250 = io_M_AXI_RDATA[127:96];
  assign _T_251 = io_M_AXI_RDATA[95:64];
  assign _T_252 = io_M_AXI_RDATA[63:32];
  assign _T_253 = io_M_AXI_RDATA[31:0];
  assign _T_279 = _T_278[5:0];
  assign _T_286 = _T_285[5:0];
  assign io_in_cmd_ready = _T_148;
  assign io_in_wdata_ready = io_M_AXI_WREADY;
  assign io_in_rresp_valid = io_M_AXI_RVALID;
  assign io_in_rresp_bits_rdata_0 = rdataAsVec_0;
  assign io_in_rresp_bits_rdata_1 = rdataAsVec_1;
  assign io_in_rresp_bits_rdata_2 = rdataAsVec_2;
  assign io_in_rresp_bits_rdata_3 = rdataAsVec_3;
  assign io_in_rresp_bits_rdata_4 = rdataAsVec_4;
  assign io_in_rresp_bits_rdata_5 = rdataAsVec_5;
  assign io_in_rresp_bits_rdata_6 = rdataAsVec_6;
  assign io_in_rresp_bits_rdata_7 = rdataAsVec_7;
  assign io_in_rresp_bits_rdata_8 = rdataAsVec_8;
  assign io_in_rresp_bits_rdata_9 = rdataAsVec_9;
  assign io_in_rresp_bits_rdata_10 = rdataAsVec_10;
  assign io_in_rresp_bits_rdata_11 = rdataAsVec_11;
  assign io_in_rresp_bits_rdata_12 = rdataAsVec_12;
  assign io_in_rresp_bits_rdata_13 = rdataAsVec_13;
  assign io_in_rresp_bits_rdata_14 = rdataAsVec_14;
  assign io_in_rresp_bits_rdata_15 = rdataAsVec_15;
  assign io_in_rresp_bits_tag_streamId = _T_276_streamId;
  assign io_in_wresp_valid = io_M_AXI_BVALID;
  assign io_in_wresp_bits_tag_streamId = _T_283_streamId;
  assign io_M_AXI_AWID = id;
  assign io_M_AXI_AWADDR = io_in_cmd_bits_addr[31:0];
  assign io_M_AXI_AWLEN = _T_139[7:0];
  assign io_M_AXI_AWVALID = _T_159;
  assign io_M_AXI_ARID = id;
  assign io_M_AXI_ARADDR = io_in_cmd_bits_addr[31:0];
  assign io_M_AXI_ARLEN = _T_139[7:0];
  assign io_M_AXI_ARVALID = _T_147;
  assign io_M_AXI_WDATA = _T_174;
  assign io_M_AXI_WSTRB = _T_237;
  assign io_M_AXI_WVALID = io_in_wdata_valid;
  assign io_M_AXI_RREADY = io_in_rresp_ready;
  assign io_M_AXI_BREADY = io_in_wresp_ready;
  assign rdataAsVec_0 = _T_253;
  assign rdataAsVec_1 = _T_252;
  assign rdataAsVec_2 = _T_251;
  assign rdataAsVec_3 = _T_250;
  assign rdataAsVec_4 = _T_249;
  assign rdataAsVec_5 = _T_248;
  assign rdataAsVec_6 = _T_247;
  assign rdataAsVec_7 = _T_246;
  assign rdataAsVec_8 = _T_245;
  assign rdataAsVec_9 = _T_244;
  assign rdataAsVec_10 = _T_243;
  assign rdataAsVec_11 = _T_242;
  assign rdataAsVec_12 = _T_241;
  assign rdataAsVec_13 = _T_240;
  assign rdataAsVec_14 = _T_239;
  assign rdataAsVec_15 = _T_238;
  assign _T_276_streamId = _T_279;
  assign _T_278 = io_M_AXI_RID;
  assign _T_283_streamId = _T_286;
  assign _T_285 = io_M_AXI_BID;
endmodule
module FringeZynq(
  input          clock,
  input          reset,
  input  [31:0]  io_S_AXI_AWADDR,
  input  [2:0]   io_S_AXI_AWPROT,
  input          io_S_AXI_AWVALID,
  output         io_S_AXI_AWREADY,
  input  [31:0]  io_S_AXI_ARADDR,
  input  [2:0]   io_S_AXI_ARPROT,
  input          io_S_AXI_ARVALID,
  output         io_S_AXI_ARREADY,
  input  [31:0]  io_S_AXI_WDATA,
  input  [3:0]   io_S_AXI_WSTRB,
  input          io_S_AXI_WVALID,
  output         io_S_AXI_WREADY,
  output [31:0]  io_S_AXI_RDATA,
  output [1:0]   io_S_AXI_RRESP,
  output         io_S_AXI_RVALID,
  input          io_S_AXI_RREADY,
  output [1:0]   io_S_AXI_BRESP,
  output         io_S_AXI_BVALID,
  input          io_S_AXI_BREADY,
  output [31:0]  io_M_AXI_0_AWID,
  output [31:0]  io_M_AXI_0_AWADDR,
  output [7:0]   io_M_AXI_0_AWLEN,
  output         io_M_AXI_0_AWVALID,
  input          io_M_AXI_0_AWREADY,
  output [31:0]  io_M_AXI_0_ARID,
  output [31:0]  io_M_AXI_0_ARADDR,
  output [7:0]   io_M_AXI_0_ARLEN,
  output         io_M_AXI_0_ARVALID,
  input          io_M_AXI_0_ARREADY,
  output [511:0] io_M_AXI_0_WDATA,
  output [63:0]  io_M_AXI_0_WSTRB,
  output         io_M_AXI_0_WVALID,
  input          io_M_AXI_0_WREADY,
  input  [31:0]  io_M_AXI_0_RID,
  input  [511:0] io_M_AXI_0_RDATA,
  input          io_M_AXI_0_RVALID,
  output         io_M_AXI_0_RREADY,
  input  [31:0]  io_M_AXI_0_BID,
  input          io_M_AXI_0_BVALID,
  output         io_M_AXI_0_BREADY,
  output [31:0]  io_M_AXI_1_AWID,
  output [31:0]  io_M_AXI_1_AWADDR,
  output [7:0]   io_M_AXI_1_AWLEN,
  output         io_M_AXI_1_AWVALID,
  input          io_M_AXI_1_AWREADY,
  output [31:0]  io_M_AXI_1_ARID,
  output [31:0]  io_M_AXI_1_ARADDR,
  output [7:0]   io_M_AXI_1_ARLEN,
  output         io_M_AXI_1_ARVALID,
  input          io_M_AXI_1_ARREADY,
  output [511:0] io_M_AXI_1_WDATA,
  output [63:0]  io_M_AXI_1_WSTRB,
  output         io_M_AXI_1_WVALID,
  input          io_M_AXI_1_WREADY,
  input  [31:0]  io_M_AXI_1_RID,
  input  [511:0] io_M_AXI_1_RDATA,
  input          io_M_AXI_1_RVALID,
  output         io_M_AXI_1_RREADY,
  input  [31:0]  io_M_AXI_1_BID,
  input          io_M_AXI_1_BVALID,
  output         io_M_AXI_1_BREADY,
  output [31:0]  io_M_AXI_2_AWID,
  output [31:0]  io_M_AXI_2_AWADDR,
  output [7:0]   io_M_AXI_2_AWLEN,
  output         io_M_AXI_2_AWVALID,
  input          io_M_AXI_2_AWREADY,
  output [31:0]  io_M_AXI_2_ARID,
  output [31:0]  io_M_AXI_2_ARADDR,
  output [7:0]   io_M_AXI_2_ARLEN,
  output         io_M_AXI_2_ARVALID,
  input          io_M_AXI_2_ARREADY,
  output [511:0] io_M_AXI_2_WDATA,
  output [63:0]  io_M_AXI_2_WSTRB,
  output         io_M_AXI_2_WVALID,
  input          io_M_AXI_2_WREADY,
  input  [31:0]  io_M_AXI_2_RID,
  input  [511:0] io_M_AXI_2_RDATA,
  input          io_M_AXI_2_RVALID,
  output         io_M_AXI_2_RREADY,
  input  [31:0]  io_M_AXI_2_BID,
  input          io_M_AXI_2_BVALID,
  output         io_M_AXI_2_BREADY,
  output [31:0]  io_M_AXI_3_AWID,
  output [31:0]  io_M_AXI_3_AWADDR,
  output [7:0]   io_M_AXI_3_AWLEN,
  output         io_M_AXI_3_AWVALID,
  input          io_M_AXI_3_AWREADY,
  output [31:0]  io_M_AXI_3_ARID,
  output [31:0]  io_M_AXI_3_ARADDR,
  output [7:0]   io_M_AXI_3_ARLEN,
  output         io_M_AXI_3_ARVALID,
  input          io_M_AXI_3_ARREADY,
  output [511:0] io_M_AXI_3_WDATA,
  output [63:0]  io_M_AXI_3_WSTRB,
  output         io_M_AXI_3_WVALID,
  input          io_M_AXI_3_WREADY,
  input  [31:0]  io_M_AXI_3_RID,
  input  [511:0] io_M_AXI_3_RDATA,
  input          io_M_AXI_3_RVALID,
  output         io_M_AXI_3_RREADY,
  input  [31:0]  io_M_AXI_3_BID,
  input          io_M_AXI_3_BVALID,
  output         io_M_AXI_3_BREADY,
  input  [31:0]  io_TOP_AXI_AWADDR,
  input  [7:0]   io_TOP_AXI_AWLEN,
  input          io_TOP_AXI_AWVALID,
  input          io_TOP_AXI_AWREADY,
  input          io_TOP_AXI_ARID,
  input  [31:0]  io_TOP_AXI_ARADDR,
  input  [7:0]   io_TOP_AXI_ARLEN,
  input  [2:0]   io_TOP_AXI_ARSIZE,
  input  [1:0]   io_TOP_AXI_ARBURST,
  input          io_TOP_AXI_ARVALID,
  input          io_TOP_AXI_ARREADY,
  input  [31:0]  io_TOP_AXI_WDATA,
  input  [63:0]  io_TOP_AXI_WSTRB,
  input          io_TOP_AXI_WVALID,
  input          io_TOP_AXI_WREADY,
  input          io_TOP_AXI_RVALID,
  input          io_TOP_AXI_RREADY,
  input          io_TOP_AXI_BVALID,
  input          io_TOP_AXI_BREADY,
  input  [31:0]  io_DWIDTH_AXI_AWADDR,
  input  [7:0]   io_DWIDTH_AXI_AWLEN,
  input          io_DWIDTH_AXI_AWVALID,
  input          io_DWIDTH_AXI_AWREADY,
  input  [31:0]  io_DWIDTH_AXI_ARADDR,
  input  [7:0]   io_DWIDTH_AXI_ARLEN,
  input  [2:0]   io_DWIDTH_AXI_ARSIZE,
  input  [1:0]   io_DWIDTH_AXI_ARBURST,
  input          io_DWIDTH_AXI_ARVALID,
  input          io_DWIDTH_AXI_ARREADY,
  input  [31:0]  io_DWIDTH_AXI_WDATA,
  input  [63:0]  io_DWIDTH_AXI_WSTRB,
  input          io_DWIDTH_AXI_WVALID,
  input          io_DWIDTH_AXI_WREADY,
  input          io_DWIDTH_AXI_RVALID,
  input          io_DWIDTH_AXI_RREADY,
  input          io_DWIDTH_AXI_BVALID,
  input          io_DWIDTH_AXI_BREADY,
  output         io_enable,
  input          io_done,
  output         io_reset,
  output [63:0]  io_argIns_0,
  output [63:0]  io_argIns_1,
  output [63:0]  io_argIns_2,
  input          io_argOuts_0_valid,
  input  [63:0]  io_argOuts_0_bits,
  output         io_memStreams_loads_3_cmd_ready,
  input          io_memStreams_loads_3_cmd_valid,
  input  [63:0]  io_memStreams_loads_3_cmd_bits_addr,
  input          io_memStreams_loads_3_cmd_bits_isWr,
  input  [15:0]  io_memStreams_loads_3_cmd_bits_size,
  input          io_memStreams_loads_3_rdata_ready,
  output         io_memStreams_loads_3_rdata_valid,
  output [31:0]  io_memStreams_loads_3_rdata_bits_0,
  output         io_memStreams_loads_2_cmd_ready,
  input          io_memStreams_loads_2_cmd_valid,
  input  [63:0]  io_memStreams_loads_2_cmd_bits_addr,
  input          io_memStreams_loads_2_cmd_bits_isWr,
  input  [15:0]  io_memStreams_loads_2_cmd_bits_size,
  input          io_memStreams_loads_2_rdata_ready,
  output         io_memStreams_loads_2_rdata_valid,
  output [31:0]  io_memStreams_loads_2_rdata_bits_0,
  output         io_memStreams_loads_1_cmd_ready,
  input          io_memStreams_loads_1_cmd_valid,
  input  [63:0]  io_memStreams_loads_1_cmd_bits_addr,
  input          io_memStreams_loads_1_cmd_bits_isWr,
  input  [15:0]  io_memStreams_loads_1_cmd_bits_size,
  input          io_memStreams_loads_1_rdata_ready,
  output         io_memStreams_loads_1_rdata_valid,
  output [31:0]  io_memStreams_loads_1_rdata_bits_0,
  output         io_memStreams_loads_0_cmd_ready,
  input          io_memStreams_loads_0_cmd_valid,
  input  [63:0]  io_memStreams_loads_0_cmd_bits_addr,
  input          io_memStreams_loads_0_cmd_bits_isWr,
  input  [15:0]  io_memStreams_loads_0_cmd_bits_size,
  input          io_memStreams_loads_0_rdata_ready,
  output         io_memStreams_loads_0_rdata_valid,
  output [31:0]  io_memStreams_loads_0_rdata_bits_0
);
  wire  fringeCommon_clock;
  wire  fringeCommon_reset;
  wire [31:0] fringeCommon_io_raddr;
  wire  fringeCommon_io_wen;
  wire [31:0] fringeCommon_io_waddr;
  wire [63:0] fringeCommon_io_wdata;
  wire [63:0] fringeCommon_io_rdata;
  wire  fringeCommon_io_enable;
  wire  fringeCommon_io_done;
  wire  fringeCommon_io_reset;
  wire [63:0] fringeCommon_io_argIns_0;
  wire [63:0] fringeCommon_io_argIns_1;
  wire [63:0] fringeCommon_io_argIns_2;
  wire  fringeCommon_io_argOuts_0_valid;
  wire [63:0] fringeCommon_io_argOuts_0_bits;
  wire  fringeCommon_io_memStreams_loads_3_cmd_ready;
  wire  fringeCommon_io_memStreams_loads_3_cmd_valid;
  wire [63:0] fringeCommon_io_memStreams_loads_3_cmd_bits_addr;
  wire  fringeCommon_io_memStreams_loads_3_cmd_bits_isWr;
  wire [15:0] fringeCommon_io_memStreams_loads_3_cmd_bits_size;
  wire  fringeCommon_io_memStreams_loads_3_rdata_ready;
  wire  fringeCommon_io_memStreams_loads_3_rdata_valid;
  wire [31:0] fringeCommon_io_memStreams_loads_3_rdata_bits_0;
  wire  fringeCommon_io_memStreams_loads_2_cmd_ready;
  wire  fringeCommon_io_memStreams_loads_2_cmd_valid;
  wire [63:0] fringeCommon_io_memStreams_loads_2_cmd_bits_addr;
  wire  fringeCommon_io_memStreams_loads_2_cmd_bits_isWr;
  wire [15:0] fringeCommon_io_memStreams_loads_2_cmd_bits_size;
  wire  fringeCommon_io_memStreams_loads_2_rdata_ready;
  wire  fringeCommon_io_memStreams_loads_2_rdata_valid;
  wire [31:0] fringeCommon_io_memStreams_loads_2_rdata_bits_0;
  wire  fringeCommon_io_memStreams_loads_1_cmd_ready;
  wire  fringeCommon_io_memStreams_loads_1_cmd_valid;
  wire [63:0] fringeCommon_io_memStreams_loads_1_cmd_bits_addr;
  wire  fringeCommon_io_memStreams_loads_1_cmd_bits_isWr;
  wire [15:0] fringeCommon_io_memStreams_loads_1_cmd_bits_size;
  wire  fringeCommon_io_memStreams_loads_1_rdata_ready;
  wire  fringeCommon_io_memStreams_loads_1_rdata_valid;
  wire [31:0] fringeCommon_io_memStreams_loads_1_rdata_bits_0;
  wire  fringeCommon_io_memStreams_loads_0_cmd_ready;
  wire  fringeCommon_io_memStreams_loads_0_cmd_valid;
  wire [63:0] fringeCommon_io_memStreams_loads_0_cmd_bits_addr;
  wire  fringeCommon_io_memStreams_loads_0_cmd_bits_isWr;
  wire [15:0] fringeCommon_io_memStreams_loads_0_cmd_bits_size;
  wire  fringeCommon_io_memStreams_loads_0_rdata_ready;
  wire  fringeCommon_io_memStreams_loads_0_rdata_valid;
  wire [31:0] fringeCommon_io_memStreams_loads_0_rdata_bits_0;
  wire  fringeCommon_io_dram_0_cmd_ready;
  wire  fringeCommon_io_dram_0_cmd_valid;
  wire [63:0] fringeCommon_io_dram_0_cmd_bits_addr;
  wire [31:0] fringeCommon_io_dram_0_cmd_bits_size;
  wire  fringeCommon_io_dram_0_cmd_bits_isWr;
  wire [25:0] fringeCommon_io_dram_0_cmd_bits_tag_uid;
  wire [5:0] fringeCommon_io_dram_0_cmd_bits_tag_streamId;
  wire  fringeCommon_io_dram_0_wdata_ready;
  wire  fringeCommon_io_dram_0_wdata_valid;
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_0;
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_1;
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_2;
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_3;
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_4;
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_5;
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_6;
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_7;
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_8;
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_9;
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_10;
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_11;
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_12;
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_13;
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_14;
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_15;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_0;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_1;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_2;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_3;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_4;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_5;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_6;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_7;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_8;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_9;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_10;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_11;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_12;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_13;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_14;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_15;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_16;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_17;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_18;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_19;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_20;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_21;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_22;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_23;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_24;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_25;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_26;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_27;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_28;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_29;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_30;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_31;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_32;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_33;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_34;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_35;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_36;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_37;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_38;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_39;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_40;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_41;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_42;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_43;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_44;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_45;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_46;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_47;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_48;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_49;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_50;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_51;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_52;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_53;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_54;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_55;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_56;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_57;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_58;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_59;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_60;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_61;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_62;
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_63;
  wire  fringeCommon_io_dram_0_rresp_ready;
  wire  fringeCommon_io_dram_0_rresp_valid;
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_rdata_0;
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_rdata_1;
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_rdata_2;
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_rdata_3;
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_rdata_4;
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_rdata_5;
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_rdata_6;
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_rdata_7;
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_rdata_8;
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_rdata_9;
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_rdata_10;
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_rdata_11;
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_rdata_12;
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_rdata_13;
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_rdata_14;
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_rdata_15;
  wire [5:0] fringeCommon_io_dram_0_rresp_bits_tag_streamId;
  wire  fringeCommon_io_dram_0_wresp_ready;
  wire  fringeCommon_io_dram_0_wresp_valid;
  wire [5:0] fringeCommon_io_dram_0_wresp_bits_tag_streamId;
  wire  fringeCommon_io_dram_1_cmd_ready;
  wire  fringeCommon_io_dram_1_cmd_valid;
  wire [63:0] fringeCommon_io_dram_1_cmd_bits_addr;
  wire [31:0] fringeCommon_io_dram_1_cmd_bits_size;
  wire  fringeCommon_io_dram_1_cmd_bits_isWr;
  wire [25:0] fringeCommon_io_dram_1_cmd_bits_tag_uid;
  wire [5:0] fringeCommon_io_dram_1_cmd_bits_tag_streamId;
  wire  fringeCommon_io_dram_1_wdata_ready;
  wire  fringeCommon_io_dram_1_wdata_valid;
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_0;
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_1;
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_2;
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_3;
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_4;
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_5;
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_6;
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_7;
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_8;
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_9;
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_10;
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_11;
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_12;
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_13;
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_14;
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_15;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_0;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_1;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_2;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_3;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_4;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_5;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_6;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_7;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_8;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_9;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_10;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_11;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_12;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_13;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_14;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_15;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_16;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_17;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_18;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_19;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_20;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_21;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_22;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_23;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_24;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_25;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_26;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_27;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_28;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_29;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_30;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_31;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_32;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_33;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_34;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_35;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_36;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_37;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_38;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_39;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_40;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_41;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_42;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_43;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_44;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_45;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_46;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_47;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_48;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_49;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_50;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_51;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_52;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_53;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_54;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_55;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_56;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_57;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_58;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_59;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_60;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_61;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_62;
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_63;
  wire  fringeCommon_io_dram_1_rresp_ready;
  wire  fringeCommon_io_dram_1_rresp_valid;
  wire [31:0] fringeCommon_io_dram_1_rresp_bits_rdata_0;
  wire [31:0] fringeCommon_io_dram_1_rresp_bits_rdata_1;
  wire [31:0] fringeCommon_io_dram_1_rresp_bits_rdata_2;
  wire [31:0] fringeCommon_io_dram_1_rresp_bits_rdata_3;
  wire [31:0] fringeCommon_io_dram_1_rresp_bits_rdata_4;
  wire [31:0] fringeCommon_io_dram_1_rresp_bits_rdata_5;
  wire [31:0] fringeCommon_io_dram_1_rresp_bits_rdata_6;
  wire [31:0] fringeCommon_io_dram_1_rresp_bits_rdata_7;
  wire [31:0] fringeCommon_io_dram_1_rresp_bits_rdata_8;
  wire [31:0] fringeCommon_io_dram_1_rresp_bits_rdata_9;
  wire [31:0] fringeCommon_io_dram_1_rresp_bits_rdata_10;
  wire [31:0] fringeCommon_io_dram_1_rresp_bits_rdata_11;
  wire [31:0] fringeCommon_io_dram_1_rresp_bits_rdata_12;
  wire [31:0] fringeCommon_io_dram_1_rresp_bits_rdata_13;
  wire [31:0] fringeCommon_io_dram_1_rresp_bits_rdata_14;
  wire [31:0] fringeCommon_io_dram_1_rresp_bits_rdata_15;
  wire [5:0] fringeCommon_io_dram_1_rresp_bits_tag_streamId;
  wire  fringeCommon_io_dram_1_wresp_ready;
  wire  fringeCommon_io_dram_1_wresp_valid;
  wire [5:0] fringeCommon_io_dram_1_wresp_bits_tag_streamId;
  wire  fringeCommon_io_dram_2_cmd_ready;
  wire  fringeCommon_io_dram_2_cmd_valid;
  wire [63:0] fringeCommon_io_dram_2_cmd_bits_addr;
  wire [31:0] fringeCommon_io_dram_2_cmd_bits_size;
  wire  fringeCommon_io_dram_2_cmd_bits_isWr;
  wire [25:0] fringeCommon_io_dram_2_cmd_bits_tag_uid;
  wire [5:0] fringeCommon_io_dram_2_cmd_bits_tag_streamId;
  wire  fringeCommon_io_dram_2_wdata_ready;
  wire  fringeCommon_io_dram_2_wdata_valid;
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_0;
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_1;
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_2;
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_3;
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_4;
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_5;
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_6;
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_7;
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_8;
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_9;
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_10;
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_11;
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_12;
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_13;
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_14;
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_15;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_0;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_1;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_2;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_3;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_4;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_5;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_6;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_7;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_8;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_9;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_10;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_11;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_12;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_13;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_14;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_15;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_16;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_17;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_18;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_19;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_20;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_21;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_22;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_23;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_24;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_25;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_26;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_27;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_28;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_29;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_30;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_31;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_32;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_33;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_34;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_35;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_36;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_37;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_38;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_39;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_40;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_41;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_42;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_43;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_44;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_45;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_46;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_47;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_48;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_49;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_50;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_51;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_52;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_53;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_54;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_55;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_56;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_57;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_58;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_59;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_60;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_61;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_62;
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_63;
  wire  fringeCommon_io_dram_2_rresp_ready;
  wire  fringeCommon_io_dram_2_rresp_valid;
  wire [31:0] fringeCommon_io_dram_2_rresp_bits_rdata_0;
  wire [31:0] fringeCommon_io_dram_2_rresp_bits_rdata_1;
  wire [31:0] fringeCommon_io_dram_2_rresp_bits_rdata_2;
  wire [31:0] fringeCommon_io_dram_2_rresp_bits_rdata_3;
  wire [31:0] fringeCommon_io_dram_2_rresp_bits_rdata_4;
  wire [31:0] fringeCommon_io_dram_2_rresp_bits_rdata_5;
  wire [31:0] fringeCommon_io_dram_2_rresp_bits_rdata_6;
  wire [31:0] fringeCommon_io_dram_2_rresp_bits_rdata_7;
  wire [31:0] fringeCommon_io_dram_2_rresp_bits_rdata_8;
  wire [31:0] fringeCommon_io_dram_2_rresp_bits_rdata_9;
  wire [31:0] fringeCommon_io_dram_2_rresp_bits_rdata_10;
  wire [31:0] fringeCommon_io_dram_2_rresp_bits_rdata_11;
  wire [31:0] fringeCommon_io_dram_2_rresp_bits_rdata_12;
  wire [31:0] fringeCommon_io_dram_2_rresp_bits_rdata_13;
  wire [31:0] fringeCommon_io_dram_2_rresp_bits_rdata_14;
  wire [31:0] fringeCommon_io_dram_2_rresp_bits_rdata_15;
  wire [5:0] fringeCommon_io_dram_2_rresp_bits_tag_streamId;
  wire  fringeCommon_io_dram_2_wresp_ready;
  wire  fringeCommon_io_dram_2_wresp_valid;
  wire [5:0] fringeCommon_io_dram_2_wresp_bits_tag_streamId;
  wire  fringeCommon_io_dram_3_cmd_ready;
  wire  fringeCommon_io_dram_3_cmd_valid;
  wire [63:0] fringeCommon_io_dram_3_cmd_bits_addr;
  wire [31:0] fringeCommon_io_dram_3_cmd_bits_size;
  wire  fringeCommon_io_dram_3_cmd_bits_isWr;
  wire [25:0] fringeCommon_io_dram_3_cmd_bits_tag_uid;
  wire [5:0] fringeCommon_io_dram_3_cmd_bits_tag_streamId;
  wire  fringeCommon_io_dram_3_wdata_ready;
  wire  fringeCommon_io_dram_3_wdata_valid;
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_0;
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_1;
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_2;
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_3;
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_4;
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_5;
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_6;
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_7;
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_8;
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_9;
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_10;
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_11;
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_12;
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_13;
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_14;
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_15;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_0;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_1;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_2;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_3;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_4;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_5;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_6;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_7;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_8;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_9;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_10;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_11;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_12;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_13;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_14;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_15;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_16;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_17;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_18;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_19;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_20;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_21;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_22;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_23;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_24;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_25;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_26;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_27;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_28;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_29;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_30;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_31;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_32;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_33;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_34;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_35;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_36;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_37;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_38;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_39;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_40;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_41;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_42;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_43;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_44;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_45;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_46;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_47;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_48;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_49;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_50;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_51;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_52;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_53;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_54;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_55;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_56;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_57;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_58;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_59;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_60;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_61;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_62;
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_63;
  wire  fringeCommon_io_dram_3_rresp_ready;
  wire  fringeCommon_io_dram_3_rresp_valid;
  wire [31:0] fringeCommon_io_dram_3_rresp_bits_rdata_0;
  wire [31:0] fringeCommon_io_dram_3_rresp_bits_rdata_1;
  wire [31:0] fringeCommon_io_dram_3_rresp_bits_rdata_2;
  wire [31:0] fringeCommon_io_dram_3_rresp_bits_rdata_3;
  wire [31:0] fringeCommon_io_dram_3_rresp_bits_rdata_4;
  wire [31:0] fringeCommon_io_dram_3_rresp_bits_rdata_5;
  wire [31:0] fringeCommon_io_dram_3_rresp_bits_rdata_6;
  wire [31:0] fringeCommon_io_dram_3_rresp_bits_rdata_7;
  wire [31:0] fringeCommon_io_dram_3_rresp_bits_rdata_8;
  wire [31:0] fringeCommon_io_dram_3_rresp_bits_rdata_9;
  wire [31:0] fringeCommon_io_dram_3_rresp_bits_rdata_10;
  wire [31:0] fringeCommon_io_dram_3_rresp_bits_rdata_11;
  wire [31:0] fringeCommon_io_dram_3_rresp_bits_rdata_12;
  wire [31:0] fringeCommon_io_dram_3_rresp_bits_rdata_13;
  wire [31:0] fringeCommon_io_dram_3_rresp_bits_rdata_14;
  wire [31:0] fringeCommon_io_dram_3_rresp_bits_rdata_15;
  wire [5:0] fringeCommon_io_dram_3_rresp_bits_tag_streamId;
  wire  fringeCommon_io_dram_3_wresp_ready;
  wire  fringeCommon_io_dram_3_wresp_valid;
  wire [5:0] fringeCommon_io_dram_3_wresp_bits_tag_streamId;
  wire [63:0] fringeCommon_io_TOP_AXI_AWADDR;
  wire [7:0] fringeCommon_io_TOP_AXI_AWLEN;
  wire  fringeCommon_io_TOP_AXI_AWVALID;
  wire  fringeCommon_io_TOP_AXI_AWREADY;
  wire  fringeCommon_io_TOP_AXI_ARID;
  wire [63:0] fringeCommon_io_TOP_AXI_ARADDR;
  wire [7:0] fringeCommon_io_TOP_AXI_ARLEN;
  wire [2:0] fringeCommon_io_TOP_AXI_ARSIZE;
  wire [1:0] fringeCommon_io_TOP_AXI_ARBURST;
  wire  fringeCommon_io_TOP_AXI_ARVALID;
  wire  fringeCommon_io_TOP_AXI_ARREADY;
  wire [511:0] fringeCommon_io_TOP_AXI_WDATA;
  wire [63:0] fringeCommon_io_TOP_AXI_WSTRB;
  wire  fringeCommon_io_TOP_AXI_WVALID;
  wire  fringeCommon_io_TOP_AXI_WREADY;
  wire  fringeCommon_io_TOP_AXI_RVALID;
  wire  fringeCommon_io_TOP_AXI_RREADY;
  wire  fringeCommon_io_TOP_AXI_BVALID;
  wire  fringeCommon_io_TOP_AXI_BREADY;
  wire [63:0] fringeCommon_io_DWIDTH_AXI_AWADDR;
  wire [7:0] fringeCommon_io_DWIDTH_AXI_AWLEN;
  wire  fringeCommon_io_DWIDTH_AXI_AWVALID;
  wire  fringeCommon_io_DWIDTH_AXI_AWREADY;
  wire [63:0] fringeCommon_io_DWIDTH_AXI_ARADDR;
  wire [7:0] fringeCommon_io_DWIDTH_AXI_ARLEN;
  wire [2:0] fringeCommon_io_DWIDTH_AXI_ARSIZE;
  wire [1:0] fringeCommon_io_DWIDTH_AXI_ARBURST;
  wire  fringeCommon_io_DWIDTH_AXI_ARVALID;
  wire  fringeCommon_io_DWIDTH_AXI_ARREADY;
  wire [511:0] fringeCommon_io_DWIDTH_AXI_WDATA;
  wire [63:0] fringeCommon_io_DWIDTH_AXI_WSTRB;
  wire  fringeCommon_io_DWIDTH_AXI_WVALID;
  wire  fringeCommon_io_DWIDTH_AXI_WREADY;
  wire  fringeCommon_io_DWIDTH_AXI_RVALID;
  wire  fringeCommon_io_DWIDTH_AXI_RREADY;
  wire  fringeCommon_io_DWIDTH_AXI_BVALID;
  wire  fringeCommon_io_DWIDTH_AXI_BREADY;
  wire  AXI4LiteToRFBridge_clock;
  wire  AXI4LiteToRFBridge_reset;
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_AWADDR;
  wire [2:0] AXI4LiteToRFBridge_io_S_AXI_AWPROT;
  wire  AXI4LiteToRFBridge_io_S_AXI_AWVALID;
  wire  AXI4LiteToRFBridge_io_S_AXI_AWREADY;
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_ARADDR;
  wire [2:0] AXI4LiteToRFBridge_io_S_AXI_ARPROT;
  wire  AXI4LiteToRFBridge_io_S_AXI_ARVALID;
  wire  AXI4LiteToRFBridge_io_S_AXI_ARREADY;
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_WDATA;
  wire [3:0] AXI4LiteToRFBridge_io_S_AXI_WSTRB;
  wire  AXI4LiteToRFBridge_io_S_AXI_WVALID;
  wire  AXI4LiteToRFBridge_io_S_AXI_WREADY;
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_RDATA;
  wire [1:0] AXI4LiteToRFBridge_io_S_AXI_RRESP;
  wire  AXI4LiteToRFBridge_io_S_AXI_RVALID;
  wire  AXI4LiteToRFBridge_io_S_AXI_RREADY;
  wire [1:0] AXI4LiteToRFBridge_io_S_AXI_BRESP;
  wire  AXI4LiteToRFBridge_io_S_AXI_BVALID;
  wire  AXI4LiteToRFBridge_io_S_AXI_BREADY;
  wire [31:0] AXI4LiteToRFBridge_io_raddr;
  wire  AXI4LiteToRFBridge_io_wen;
  wire [31:0] AXI4LiteToRFBridge_io_waddr;
  wire [31:0] AXI4LiteToRFBridge_io_wdata;
  wire [31:0] AXI4LiteToRFBridge_io_rdata;
  wire  MAGToAXI4Bridge_io_in_cmd_ready;
  wire  MAGToAXI4Bridge_io_in_cmd_valid;
  wire [63:0] MAGToAXI4Bridge_io_in_cmd_bits_addr;
  wire [31:0] MAGToAXI4Bridge_io_in_cmd_bits_size;
  wire  MAGToAXI4Bridge_io_in_cmd_bits_isWr;
  wire [25:0] MAGToAXI4Bridge_io_in_cmd_bits_tag_uid;
  wire [5:0] MAGToAXI4Bridge_io_in_cmd_bits_tag_streamId;
  wire  MAGToAXI4Bridge_io_in_wdata_ready;
  wire  MAGToAXI4Bridge_io_in_wdata_valid;
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_0;
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_1;
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_2;
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_3;
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_4;
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_5;
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_6;
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_7;
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_8;
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_9;
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_10;
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_11;
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_12;
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_13;
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_14;
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_15;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_0;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_1;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_2;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_3;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_4;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_5;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_6;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_7;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_8;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_9;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_10;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_11;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_12;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_13;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_14;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_15;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_16;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_17;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_18;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_19;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_20;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_21;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_22;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_23;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_24;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_25;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_26;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_27;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_28;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_29;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_30;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_31;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_32;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_33;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_34;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_35;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_36;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_37;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_38;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_39;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_40;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_41;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_42;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_43;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_44;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_45;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_46;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_47;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_48;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_49;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_50;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_51;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_52;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_53;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_54;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_55;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_56;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_57;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_58;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_59;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_60;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_61;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_62;
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_63;
  wire  MAGToAXI4Bridge_io_in_rresp_ready;
  wire  MAGToAXI4Bridge_io_in_rresp_valid;
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_0;
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_1;
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_2;
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_3;
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_4;
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_5;
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_6;
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_7;
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_8;
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_9;
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_10;
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_11;
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_12;
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_13;
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_14;
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_15;
  wire [5:0] MAGToAXI4Bridge_io_in_rresp_bits_tag_streamId;
  wire  MAGToAXI4Bridge_io_in_wresp_ready;
  wire  MAGToAXI4Bridge_io_in_wresp_valid;
  wire [5:0] MAGToAXI4Bridge_io_in_wresp_bits_tag_streamId;
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_AWID;
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_AWADDR;
  wire [7:0] MAGToAXI4Bridge_io_M_AXI_AWLEN;
  wire  MAGToAXI4Bridge_io_M_AXI_AWVALID;
  wire  MAGToAXI4Bridge_io_M_AXI_AWREADY;
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_ARID;
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_ARADDR;
  wire [7:0] MAGToAXI4Bridge_io_M_AXI_ARLEN;
  wire  MAGToAXI4Bridge_io_M_AXI_ARVALID;
  wire  MAGToAXI4Bridge_io_M_AXI_ARREADY;
  wire [511:0] MAGToAXI4Bridge_io_M_AXI_WDATA;
  wire [63:0] MAGToAXI4Bridge_io_M_AXI_WSTRB;
  wire  MAGToAXI4Bridge_io_M_AXI_WVALID;
  wire  MAGToAXI4Bridge_io_M_AXI_WREADY;
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_RID;
  wire [511:0] MAGToAXI4Bridge_io_M_AXI_RDATA;
  wire  MAGToAXI4Bridge_io_M_AXI_RVALID;
  wire  MAGToAXI4Bridge_io_M_AXI_RREADY;
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_BID;
  wire  MAGToAXI4Bridge_io_M_AXI_BVALID;
  wire  MAGToAXI4Bridge_io_M_AXI_BREADY;
  wire  MAGToAXI4Bridge_1_io_in_cmd_ready;
  wire  MAGToAXI4Bridge_1_io_in_cmd_valid;
  wire [63:0] MAGToAXI4Bridge_1_io_in_cmd_bits_addr;
  wire [31:0] MAGToAXI4Bridge_1_io_in_cmd_bits_size;
  wire  MAGToAXI4Bridge_1_io_in_cmd_bits_isWr;
  wire [25:0] MAGToAXI4Bridge_1_io_in_cmd_bits_tag_uid;
  wire [5:0] MAGToAXI4Bridge_1_io_in_cmd_bits_tag_streamId;
  wire  MAGToAXI4Bridge_1_io_in_wdata_ready;
  wire  MAGToAXI4Bridge_1_io_in_wdata_valid;
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_0;
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_1;
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_2;
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_3;
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_4;
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_5;
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_6;
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_7;
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_8;
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_9;
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_10;
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_11;
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_12;
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_13;
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_14;
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_15;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_0;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_1;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_2;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_3;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_4;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_5;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_6;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_7;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_8;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_9;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_10;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_11;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_12;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_13;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_14;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_15;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_16;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_17;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_18;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_19;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_20;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_21;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_22;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_23;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_24;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_25;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_26;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_27;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_28;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_29;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_30;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_31;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_32;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_33;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_34;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_35;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_36;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_37;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_38;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_39;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_40;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_41;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_42;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_43;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_44;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_45;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_46;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_47;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_48;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_49;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_50;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_51;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_52;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_53;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_54;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_55;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_56;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_57;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_58;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_59;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_60;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_61;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_62;
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_63;
  wire  MAGToAXI4Bridge_1_io_in_rresp_ready;
  wire  MAGToAXI4Bridge_1_io_in_rresp_valid;
  wire [31:0] MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_0;
  wire [31:0] MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_1;
  wire [31:0] MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_2;
  wire [31:0] MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_3;
  wire [31:0] MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_4;
  wire [31:0] MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_5;
  wire [31:0] MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_6;
  wire [31:0] MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_7;
  wire [31:0] MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_8;
  wire [31:0] MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_9;
  wire [31:0] MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_10;
  wire [31:0] MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_11;
  wire [31:0] MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_12;
  wire [31:0] MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_13;
  wire [31:0] MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_14;
  wire [31:0] MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_15;
  wire [5:0] MAGToAXI4Bridge_1_io_in_rresp_bits_tag_streamId;
  wire  MAGToAXI4Bridge_1_io_in_wresp_ready;
  wire  MAGToAXI4Bridge_1_io_in_wresp_valid;
  wire [5:0] MAGToAXI4Bridge_1_io_in_wresp_bits_tag_streamId;
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_AWID;
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_AWADDR;
  wire [7:0] MAGToAXI4Bridge_1_io_M_AXI_AWLEN;
  wire  MAGToAXI4Bridge_1_io_M_AXI_AWVALID;
  wire  MAGToAXI4Bridge_1_io_M_AXI_AWREADY;
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_ARID;
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_ARADDR;
  wire [7:0] MAGToAXI4Bridge_1_io_M_AXI_ARLEN;
  wire  MAGToAXI4Bridge_1_io_M_AXI_ARVALID;
  wire  MAGToAXI4Bridge_1_io_M_AXI_ARREADY;
  wire [511:0] MAGToAXI4Bridge_1_io_M_AXI_WDATA;
  wire [63:0] MAGToAXI4Bridge_1_io_M_AXI_WSTRB;
  wire  MAGToAXI4Bridge_1_io_M_AXI_WVALID;
  wire  MAGToAXI4Bridge_1_io_M_AXI_WREADY;
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_RID;
  wire [511:0] MAGToAXI4Bridge_1_io_M_AXI_RDATA;
  wire  MAGToAXI4Bridge_1_io_M_AXI_RVALID;
  wire  MAGToAXI4Bridge_1_io_M_AXI_RREADY;
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_BID;
  wire  MAGToAXI4Bridge_1_io_M_AXI_BVALID;
  wire  MAGToAXI4Bridge_1_io_M_AXI_BREADY;
  wire  MAGToAXI4Bridge_2_io_in_cmd_ready;
  wire  MAGToAXI4Bridge_2_io_in_cmd_valid;
  wire [63:0] MAGToAXI4Bridge_2_io_in_cmd_bits_addr;
  wire [31:0] MAGToAXI4Bridge_2_io_in_cmd_bits_size;
  wire  MAGToAXI4Bridge_2_io_in_cmd_bits_isWr;
  wire [25:0] MAGToAXI4Bridge_2_io_in_cmd_bits_tag_uid;
  wire [5:0] MAGToAXI4Bridge_2_io_in_cmd_bits_tag_streamId;
  wire  MAGToAXI4Bridge_2_io_in_wdata_ready;
  wire  MAGToAXI4Bridge_2_io_in_wdata_valid;
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_0;
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_1;
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_2;
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_3;
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_4;
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_5;
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_6;
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_7;
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_8;
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_9;
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_10;
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_11;
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_12;
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_13;
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_14;
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_15;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_0;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_1;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_2;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_3;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_4;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_5;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_6;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_7;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_8;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_9;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_10;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_11;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_12;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_13;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_14;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_15;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_16;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_17;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_18;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_19;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_20;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_21;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_22;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_23;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_24;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_25;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_26;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_27;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_28;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_29;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_30;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_31;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_32;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_33;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_34;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_35;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_36;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_37;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_38;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_39;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_40;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_41;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_42;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_43;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_44;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_45;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_46;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_47;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_48;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_49;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_50;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_51;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_52;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_53;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_54;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_55;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_56;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_57;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_58;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_59;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_60;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_61;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_62;
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_63;
  wire  MAGToAXI4Bridge_2_io_in_rresp_ready;
  wire  MAGToAXI4Bridge_2_io_in_rresp_valid;
  wire [31:0] MAGToAXI4Bridge_2_io_in_rresp_bits_rdata_0;
  wire [31:0] MAGToAXI4Bridge_2_io_in_rresp_bits_rdata_1;
  wire [31:0] MAGToAXI4Bridge_2_io_in_rresp_bits_rdata_2;
  wire [31:0] MAGToAXI4Bridge_2_io_in_rresp_bits_rdata_3;
  wire [31:0] MAGToAXI4Bridge_2_io_in_rresp_bits_rdata_4;
  wire [31:0] MAGToAXI4Bridge_2_io_in_rresp_bits_rdata_5;
  wire [31:0] MAGToAXI4Bridge_2_io_in_rresp_bits_rdata_6;
  wire [31:0] MAGToAXI4Bridge_2_io_in_rresp_bits_rdata_7;
  wire [31:0] MAGToAXI4Bridge_2_io_in_rresp_bits_rdata_8;
  wire [31:0] MAGToAXI4Bridge_2_io_in_rresp_bits_rdata_9;
  wire [31:0] MAGToAXI4Bridge_2_io_in_rresp_bits_rdata_10;
  wire [31:0] MAGToAXI4Bridge_2_io_in_rresp_bits_rdata_11;
  wire [31:0] MAGToAXI4Bridge_2_io_in_rresp_bits_rdata_12;
  wire [31:0] MAGToAXI4Bridge_2_io_in_rresp_bits_rdata_13;
  wire [31:0] MAGToAXI4Bridge_2_io_in_rresp_bits_rdata_14;
  wire [31:0] MAGToAXI4Bridge_2_io_in_rresp_bits_rdata_15;
  wire [5:0] MAGToAXI4Bridge_2_io_in_rresp_bits_tag_streamId;
  wire  MAGToAXI4Bridge_2_io_in_wresp_ready;
  wire  MAGToAXI4Bridge_2_io_in_wresp_valid;
  wire [5:0] MAGToAXI4Bridge_2_io_in_wresp_bits_tag_streamId;
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_AWID;
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_AWADDR;
  wire [7:0] MAGToAXI4Bridge_2_io_M_AXI_AWLEN;
  wire  MAGToAXI4Bridge_2_io_M_AXI_AWVALID;
  wire  MAGToAXI4Bridge_2_io_M_AXI_AWREADY;
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_ARID;
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_ARADDR;
  wire [7:0] MAGToAXI4Bridge_2_io_M_AXI_ARLEN;
  wire  MAGToAXI4Bridge_2_io_M_AXI_ARVALID;
  wire  MAGToAXI4Bridge_2_io_M_AXI_ARREADY;
  wire [511:0] MAGToAXI4Bridge_2_io_M_AXI_WDATA;
  wire [63:0] MAGToAXI4Bridge_2_io_M_AXI_WSTRB;
  wire  MAGToAXI4Bridge_2_io_M_AXI_WVALID;
  wire  MAGToAXI4Bridge_2_io_M_AXI_WREADY;
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_RID;
  wire [511:0] MAGToAXI4Bridge_2_io_M_AXI_RDATA;
  wire  MAGToAXI4Bridge_2_io_M_AXI_RVALID;
  wire  MAGToAXI4Bridge_2_io_M_AXI_RREADY;
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_BID;
  wire  MAGToAXI4Bridge_2_io_M_AXI_BVALID;
  wire  MAGToAXI4Bridge_2_io_M_AXI_BREADY;
  wire  MAGToAXI4Bridge_3_io_in_cmd_ready;
  wire  MAGToAXI4Bridge_3_io_in_cmd_valid;
  wire [63:0] MAGToAXI4Bridge_3_io_in_cmd_bits_addr;
  wire [31:0] MAGToAXI4Bridge_3_io_in_cmd_bits_size;
  wire  MAGToAXI4Bridge_3_io_in_cmd_bits_isWr;
  wire [25:0] MAGToAXI4Bridge_3_io_in_cmd_bits_tag_uid;
  wire [5:0] MAGToAXI4Bridge_3_io_in_cmd_bits_tag_streamId;
  wire  MAGToAXI4Bridge_3_io_in_wdata_ready;
  wire  MAGToAXI4Bridge_3_io_in_wdata_valid;
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_0;
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_1;
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_2;
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_3;
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_4;
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_5;
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_6;
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_7;
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_8;
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_9;
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_10;
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_11;
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_12;
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_13;
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_14;
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_15;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_0;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_1;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_2;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_3;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_4;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_5;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_6;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_7;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_8;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_9;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_10;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_11;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_12;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_13;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_14;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_15;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_16;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_17;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_18;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_19;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_20;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_21;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_22;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_23;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_24;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_25;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_26;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_27;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_28;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_29;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_30;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_31;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_32;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_33;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_34;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_35;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_36;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_37;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_38;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_39;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_40;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_41;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_42;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_43;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_44;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_45;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_46;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_47;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_48;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_49;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_50;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_51;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_52;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_53;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_54;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_55;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_56;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_57;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_58;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_59;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_60;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_61;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_62;
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_63;
  wire  MAGToAXI4Bridge_3_io_in_rresp_ready;
  wire  MAGToAXI4Bridge_3_io_in_rresp_valid;
  wire [31:0] MAGToAXI4Bridge_3_io_in_rresp_bits_rdata_0;
  wire [31:0] MAGToAXI4Bridge_3_io_in_rresp_bits_rdata_1;
  wire [31:0] MAGToAXI4Bridge_3_io_in_rresp_bits_rdata_2;
  wire [31:0] MAGToAXI4Bridge_3_io_in_rresp_bits_rdata_3;
  wire [31:0] MAGToAXI4Bridge_3_io_in_rresp_bits_rdata_4;
  wire [31:0] MAGToAXI4Bridge_3_io_in_rresp_bits_rdata_5;
  wire [31:0] MAGToAXI4Bridge_3_io_in_rresp_bits_rdata_6;
  wire [31:0] MAGToAXI4Bridge_3_io_in_rresp_bits_rdata_7;
  wire [31:0] MAGToAXI4Bridge_3_io_in_rresp_bits_rdata_8;
  wire [31:0] MAGToAXI4Bridge_3_io_in_rresp_bits_rdata_9;
  wire [31:0] MAGToAXI4Bridge_3_io_in_rresp_bits_rdata_10;
  wire [31:0] MAGToAXI4Bridge_3_io_in_rresp_bits_rdata_11;
  wire [31:0] MAGToAXI4Bridge_3_io_in_rresp_bits_rdata_12;
  wire [31:0] MAGToAXI4Bridge_3_io_in_rresp_bits_rdata_13;
  wire [31:0] MAGToAXI4Bridge_3_io_in_rresp_bits_rdata_14;
  wire [31:0] MAGToAXI4Bridge_3_io_in_rresp_bits_rdata_15;
  wire [5:0] MAGToAXI4Bridge_3_io_in_rresp_bits_tag_streamId;
  wire  MAGToAXI4Bridge_3_io_in_wresp_ready;
  wire  MAGToAXI4Bridge_3_io_in_wresp_valid;
  wire [5:0] MAGToAXI4Bridge_3_io_in_wresp_bits_tag_streamId;
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_AWID;
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_AWADDR;
  wire [7:0] MAGToAXI4Bridge_3_io_M_AXI_AWLEN;
  wire  MAGToAXI4Bridge_3_io_M_AXI_AWVALID;
  wire  MAGToAXI4Bridge_3_io_M_AXI_AWREADY;
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_ARID;
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_ARADDR;
  wire [7:0] MAGToAXI4Bridge_3_io_M_AXI_ARLEN;
  wire  MAGToAXI4Bridge_3_io_M_AXI_ARVALID;
  wire  MAGToAXI4Bridge_3_io_M_AXI_ARREADY;
  wire [511:0] MAGToAXI4Bridge_3_io_M_AXI_WDATA;
  wire [63:0] MAGToAXI4Bridge_3_io_M_AXI_WSTRB;
  wire  MAGToAXI4Bridge_3_io_M_AXI_WVALID;
  wire  MAGToAXI4Bridge_3_io_M_AXI_WREADY;
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_RID;
  wire [511:0] MAGToAXI4Bridge_3_io_M_AXI_RDATA;
  wire  MAGToAXI4Bridge_3_io_M_AXI_RVALID;
  wire  MAGToAXI4Bridge_3_io_M_AXI_RREADY;
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_BID;
  wire  MAGToAXI4Bridge_3_io_M_AXI_BVALID;
  wire  MAGToAXI4Bridge_3_io_M_AXI_BREADY;
  Fringe fringeCommon (
    .clock(fringeCommon_clock),
    .reset(fringeCommon_reset),
    .io_raddr(fringeCommon_io_raddr),
    .io_wen(fringeCommon_io_wen),
    .io_waddr(fringeCommon_io_waddr),
    .io_wdata(fringeCommon_io_wdata),
    .io_rdata(fringeCommon_io_rdata),
    .io_enable(fringeCommon_io_enable),
    .io_done(fringeCommon_io_done),
    .io_reset(fringeCommon_io_reset),
    .io_argIns_0(fringeCommon_io_argIns_0),
    .io_argIns_1(fringeCommon_io_argIns_1),
    .io_argIns_2(fringeCommon_io_argIns_2),
    .io_argOuts_0_valid(fringeCommon_io_argOuts_0_valid),
    .io_argOuts_0_bits(fringeCommon_io_argOuts_0_bits),
    .io_memStreams_loads_3_cmd_ready(fringeCommon_io_memStreams_loads_3_cmd_ready),
    .io_memStreams_loads_3_cmd_valid(fringeCommon_io_memStreams_loads_3_cmd_valid),
    .io_memStreams_loads_3_cmd_bits_addr(fringeCommon_io_memStreams_loads_3_cmd_bits_addr),
    .io_memStreams_loads_3_cmd_bits_isWr(fringeCommon_io_memStreams_loads_3_cmd_bits_isWr),
    .io_memStreams_loads_3_cmd_bits_size(fringeCommon_io_memStreams_loads_3_cmd_bits_size),
    .io_memStreams_loads_3_rdata_ready(fringeCommon_io_memStreams_loads_3_rdata_ready),
    .io_memStreams_loads_3_rdata_valid(fringeCommon_io_memStreams_loads_3_rdata_valid),
    .io_memStreams_loads_3_rdata_bits_0(fringeCommon_io_memStreams_loads_3_rdata_bits_0),
    .io_memStreams_loads_2_cmd_ready(fringeCommon_io_memStreams_loads_2_cmd_ready),
    .io_memStreams_loads_2_cmd_valid(fringeCommon_io_memStreams_loads_2_cmd_valid),
    .io_memStreams_loads_2_cmd_bits_addr(fringeCommon_io_memStreams_loads_2_cmd_bits_addr),
    .io_memStreams_loads_2_cmd_bits_isWr(fringeCommon_io_memStreams_loads_2_cmd_bits_isWr),
    .io_memStreams_loads_2_cmd_bits_size(fringeCommon_io_memStreams_loads_2_cmd_bits_size),
    .io_memStreams_loads_2_rdata_ready(fringeCommon_io_memStreams_loads_2_rdata_ready),
    .io_memStreams_loads_2_rdata_valid(fringeCommon_io_memStreams_loads_2_rdata_valid),
    .io_memStreams_loads_2_rdata_bits_0(fringeCommon_io_memStreams_loads_2_rdata_bits_0),
    .io_memStreams_loads_1_cmd_ready(fringeCommon_io_memStreams_loads_1_cmd_ready),
    .io_memStreams_loads_1_cmd_valid(fringeCommon_io_memStreams_loads_1_cmd_valid),
    .io_memStreams_loads_1_cmd_bits_addr(fringeCommon_io_memStreams_loads_1_cmd_bits_addr),
    .io_memStreams_loads_1_cmd_bits_isWr(fringeCommon_io_memStreams_loads_1_cmd_bits_isWr),
    .io_memStreams_loads_1_cmd_bits_size(fringeCommon_io_memStreams_loads_1_cmd_bits_size),
    .io_memStreams_loads_1_rdata_ready(fringeCommon_io_memStreams_loads_1_rdata_ready),
    .io_memStreams_loads_1_rdata_valid(fringeCommon_io_memStreams_loads_1_rdata_valid),
    .io_memStreams_loads_1_rdata_bits_0(fringeCommon_io_memStreams_loads_1_rdata_bits_0),
    .io_memStreams_loads_0_cmd_ready(fringeCommon_io_memStreams_loads_0_cmd_ready),
    .io_memStreams_loads_0_cmd_valid(fringeCommon_io_memStreams_loads_0_cmd_valid),
    .io_memStreams_loads_0_cmd_bits_addr(fringeCommon_io_memStreams_loads_0_cmd_bits_addr),
    .io_memStreams_loads_0_cmd_bits_isWr(fringeCommon_io_memStreams_loads_0_cmd_bits_isWr),
    .io_memStreams_loads_0_cmd_bits_size(fringeCommon_io_memStreams_loads_0_cmd_bits_size),
    .io_memStreams_loads_0_rdata_ready(fringeCommon_io_memStreams_loads_0_rdata_ready),
    .io_memStreams_loads_0_rdata_valid(fringeCommon_io_memStreams_loads_0_rdata_valid),
    .io_memStreams_loads_0_rdata_bits_0(fringeCommon_io_memStreams_loads_0_rdata_bits_0),
    .io_dram_0_cmd_ready(fringeCommon_io_dram_0_cmd_ready),
    .io_dram_0_cmd_valid(fringeCommon_io_dram_0_cmd_valid),
    .io_dram_0_cmd_bits_addr(fringeCommon_io_dram_0_cmd_bits_addr),
    .io_dram_0_cmd_bits_size(fringeCommon_io_dram_0_cmd_bits_size),
    .io_dram_0_cmd_bits_isWr(fringeCommon_io_dram_0_cmd_bits_isWr),
    .io_dram_0_cmd_bits_tag_uid(fringeCommon_io_dram_0_cmd_bits_tag_uid),
    .io_dram_0_cmd_bits_tag_streamId(fringeCommon_io_dram_0_cmd_bits_tag_streamId),
    .io_dram_0_wdata_ready(fringeCommon_io_dram_0_wdata_ready),
    .io_dram_0_wdata_valid(fringeCommon_io_dram_0_wdata_valid),
    .io_dram_0_wdata_bits_wdata_0(fringeCommon_io_dram_0_wdata_bits_wdata_0),
    .io_dram_0_wdata_bits_wdata_1(fringeCommon_io_dram_0_wdata_bits_wdata_1),
    .io_dram_0_wdata_bits_wdata_2(fringeCommon_io_dram_0_wdata_bits_wdata_2),
    .io_dram_0_wdata_bits_wdata_3(fringeCommon_io_dram_0_wdata_bits_wdata_3),
    .io_dram_0_wdata_bits_wdata_4(fringeCommon_io_dram_0_wdata_bits_wdata_4),
    .io_dram_0_wdata_bits_wdata_5(fringeCommon_io_dram_0_wdata_bits_wdata_5),
    .io_dram_0_wdata_bits_wdata_6(fringeCommon_io_dram_0_wdata_bits_wdata_6),
    .io_dram_0_wdata_bits_wdata_7(fringeCommon_io_dram_0_wdata_bits_wdata_7),
    .io_dram_0_wdata_bits_wdata_8(fringeCommon_io_dram_0_wdata_bits_wdata_8),
    .io_dram_0_wdata_bits_wdata_9(fringeCommon_io_dram_0_wdata_bits_wdata_9),
    .io_dram_0_wdata_bits_wdata_10(fringeCommon_io_dram_0_wdata_bits_wdata_10),
    .io_dram_0_wdata_bits_wdata_11(fringeCommon_io_dram_0_wdata_bits_wdata_11),
    .io_dram_0_wdata_bits_wdata_12(fringeCommon_io_dram_0_wdata_bits_wdata_12),
    .io_dram_0_wdata_bits_wdata_13(fringeCommon_io_dram_0_wdata_bits_wdata_13),
    .io_dram_0_wdata_bits_wdata_14(fringeCommon_io_dram_0_wdata_bits_wdata_14),
    .io_dram_0_wdata_bits_wdata_15(fringeCommon_io_dram_0_wdata_bits_wdata_15),
    .io_dram_0_wdata_bits_wstrb_0(fringeCommon_io_dram_0_wdata_bits_wstrb_0),
    .io_dram_0_wdata_bits_wstrb_1(fringeCommon_io_dram_0_wdata_bits_wstrb_1),
    .io_dram_0_wdata_bits_wstrb_2(fringeCommon_io_dram_0_wdata_bits_wstrb_2),
    .io_dram_0_wdata_bits_wstrb_3(fringeCommon_io_dram_0_wdata_bits_wstrb_3),
    .io_dram_0_wdata_bits_wstrb_4(fringeCommon_io_dram_0_wdata_bits_wstrb_4),
    .io_dram_0_wdata_bits_wstrb_5(fringeCommon_io_dram_0_wdata_bits_wstrb_5),
    .io_dram_0_wdata_bits_wstrb_6(fringeCommon_io_dram_0_wdata_bits_wstrb_6),
    .io_dram_0_wdata_bits_wstrb_7(fringeCommon_io_dram_0_wdata_bits_wstrb_7),
    .io_dram_0_wdata_bits_wstrb_8(fringeCommon_io_dram_0_wdata_bits_wstrb_8),
    .io_dram_0_wdata_bits_wstrb_9(fringeCommon_io_dram_0_wdata_bits_wstrb_9),
    .io_dram_0_wdata_bits_wstrb_10(fringeCommon_io_dram_0_wdata_bits_wstrb_10),
    .io_dram_0_wdata_bits_wstrb_11(fringeCommon_io_dram_0_wdata_bits_wstrb_11),
    .io_dram_0_wdata_bits_wstrb_12(fringeCommon_io_dram_0_wdata_bits_wstrb_12),
    .io_dram_0_wdata_bits_wstrb_13(fringeCommon_io_dram_0_wdata_bits_wstrb_13),
    .io_dram_0_wdata_bits_wstrb_14(fringeCommon_io_dram_0_wdata_bits_wstrb_14),
    .io_dram_0_wdata_bits_wstrb_15(fringeCommon_io_dram_0_wdata_bits_wstrb_15),
    .io_dram_0_wdata_bits_wstrb_16(fringeCommon_io_dram_0_wdata_bits_wstrb_16),
    .io_dram_0_wdata_bits_wstrb_17(fringeCommon_io_dram_0_wdata_bits_wstrb_17),
    .io_dram_0_wdata_bits_wstrb_18(fringeCommon_io_dram_0_wdata_bits_wstrb_18),
    .io_dram_0_wdata_bits_wstrb_19(fringeCommon_io_dram_0_wdata_bits_wstrb_19),
    .io_dram_0_wdata_bits_wstrb_20(fringeCommon_io_dram_0_wdata_bits_wstrb_20),
    .io_dram_0_wdata_bits_wstrb_21(fringeCommon_io_dram_0_wdata_bits_wstrb_21),
    .io_dram_0_wdata_bits_wstrb_22(fringeCommon_io_dram_0_wdata_bits_wstrb_22),
    .io_dram_0_wdata_bits_wstrb_23(fringeCommon_io_dram_0_wdata_bits_wstrb_23),
    .io_dram_0_wdata_bits_wstrb_24(fringeCommon_io_dram_0_wdata_bits_wstrb_24),
    .io_dram_0_wdata_bits_wstrb_25(fringeCommon_io_dram_0_wdata_bits_wstrb_25),
    .io_dram_0_wdata_bits_wstrb_26(fringeCommon_io_dram_0_wdata_bits_wstrb_26),
    .io_dram_0_wdata_bits_wstrb_27(fringeCommon_io_dram_0_wdata_bits_wstrb_27),
    .io_dram_0_wdata_bits_wstrb_28(fringeCommon_io_dram_0_wdata_bits_wstrb_28),
    .io_dram_0_wdata_bits_wstrb_29(fringeCommon_io_dram_0_wdata_bits_wstrb_29),
    .io_dram_0_wdata_bits_wstrb_30(fringeCommon_io_dram_0_wdata_bits_wstrb_30),
    .io_dram_0_wdata_bits_wstrb_31(fringeCommon_io_dram_0_wdata_bits_wstrb_31),
    .io_dram_0_wdata_bits_wstrb_32(fringeCommon_io_dram_0_wdata_bits_wstrb_32),
    .io_dram_0_wdata_bits_wstrb_33(fringeCommon_io_dram_0_wdata_bits_wstrb_33),
    .io_dram_0_wdata_bits_wstrb_34(fringeCommon_io_dram_0_wdata_bits_wstrb_34),
    .io_dram_0_wdata_bits_wstrb_35(fringeCommon_io_dram_0_wdata_bits_wstrb_35),
    .io_dram_0_wdata_bits_wstrb_36(fringeCommon_io_dram_0_wdata_bits_wstrb_36),
    .io_dram_0_wdata_bits_wstrb_37(fringeCommon_io_dram_0_wdata_bits_wstrb_37),
    .io_dram_0_wdata_bits_wstrb_38(fringeCommon_io_dram_0_wdata_bits_wstrb_38),
    .io_dram_0_wdata_bits_wstrb_39(fringeCommon_io_dram_0_wdata_bits_wstrb_39),
    .io_dram_0_wdata_bits_wstrb_40(fringeCommon_io_dram_0_wdata_bits_wstrb_40),
    .io_dram_0_wdata_bits_wstrb_41(fringeCommon_io_dram_0_wdata_bits_wstrb_41),
    .io_dram_0_wdata_bits_wstrb_42(fringeCommon_io_dram_0_wdata_bits_wstrb_42),
    .io_dram_0_wdata_bits_wstrb_43(fringeCommon_io_dram_0_wdata_bits_wstrb_43),
    .io_dram_0_wdata_bits_wstrb_44(fringeCommon_io_dram_0_wdata_bits_wstrb_44),
    .io_dram_0_wdata_bits_wstrb_45(fringeCommon_io_dram_0_wdata_bits_wstrb_45),
    .io_dram_0_wdata_bits_wstrb_46(fringeCommon_io_dram_0_wdata_bits_wstrb_46),
    .io_dram_0_wdata_bits_wstrb_47(fringeCommon_io_dram_0_wdata_bits_wstrb_47),
    .io_dram_0_wdata_bits_wstrb_48(fringeCommon_io_dram_0_wdata_bits_wstrb_48),
    .io_dram_0_wdata_bits_wstrb_49(fringeCommon_io_dram_0_wdata_bits_wstrb_49),
    .io_dram_0_wdata_bits_wstrb_50(fringeCommon_io_dram_0_wdata_bits_wstrb_50),
    .io_dram_0_wdata_bits_wstrb_51(fringeCommon_io_dram_0_wdata_bits_wstrb_51),
    .io_dram_0_wdata_bits_wstrb_52(fringeCommon_io_dram_0_wdata_bits_wstrb_52),
    .io_dram_0_wdata_bits_wstrb_53(fringeCommon_io_dram_0_wdata_bits_wstrb_53),
    .io_dram_0_wdata_bits_wstrb_54(fringeCommon_io_dram_0_wdata_bits_wstrb_54),
    .io_dram_0_wdata_bits_wstrb_55(fringeCommon_io_dram_0_wdata_bits_wstrb_55),
    .io_dram_0_wdata_bits_wstrb_56(fringeCommon_io_dram_0_wdata_bits_wstrb_56),
    .io_dram_0_wdata_bits_wstrb_57(fringeCommon_io_dram_0_wdata_bits_wstrb_57),
    .io_dram_0_wdata_bits_wstrb_58(fringeCommon_io_dram_0_wdata_bits_wstrb_58),
    .io_dram_0_wdata_bits_wstrb_59(fringeCommon_io_dram_0_wdata_bits_wstrb_59),
    .io_dram_0_wdata_bits_wstrb_60(fringeCommon_io_dram_0_wdata_bits_wstrb_60),
    .io_dram_0_wdata_bits_wstrb_61(fringeCommon_io_dram_0_wdata_bits_wstrb_61),
    .io_dram_0_wdata_bits_wstrb_62(fringeCommon_io_dram_0_wdata_bits_wstrb_62),
    .io_dram_0_wdata_bits_wstrb_63(fringeCommon_io_dram_0_wdata_bits_wstrb_63),
    .io_dram_0_rresp_ready(fringeCommon_io_dram_0_rresp_ready),
    .io_dram_0_rresp_valid(fringeCommon_io_dram_0_rresp_valid),
    .io_dram_0_rresp_bits_rdata_0(fringeCommon_io_dram_0_rresp_bits_rdata_0),
    .io_dram_0_rresp_bits_rdata_1(fringeCommon_io_dram_0_rresp_bits_rdata_1),
    .io_dram_0_rresp_bits_rdata_2(fringeCommon_io_dram_0_rresp_bits_rdata_2),
    .io_dram_0_rresp_bits_rdata_3(fringeCommon_io_dram_0_rresp_bits_rdata_3),
    .io_dram_0_rresp_bits_rdata_4(fringeCommon_io_dram_0_rresp_bits_rdata_4),
    .io_dram_0_rresp_bits_rdata_5(fringeCommon_io_dram_0_rresp_bits_rdata_5),
    .io_dram_0_rresp_bits_rdata_6(fringeCommon_io_dram_0_rresp_bits_rdata_6),
    .io_dram_0_rresp_bits_rdata_7(fringeCommon_io_dram_0_rresp_bits_rdata_7),
    .io_dram_0_rresp_bits_rdata_8(fringeCommon_io_dram_0_rresp_bits_rdata_8),
    .io_dram_0_rresp_bits_rdata_9(fringeCommon_io_dram_0_rresp_bits_rdata_9),
    .io_dram_0_rresp_bits_rdata_10(fringeCommon_io_dram_0_rresp_bits_rdata_10),
    .io_dram_0_rresp_bits_rdata_11(fringeCommon_io_dram_0_rresp_bits_rdata_11),
    .io_dram_0_rresp_bits_rdata_12(fringeCommon_io_dram_0_rresp_bits_rdata_12),
    .io_dram_0_rresp_bits_rdata_13(fringeCommon_io_dram_0_rresp_bits_rdata_13),
    .io_dram_0_rresp_bits_rdata_14(fringeCommon_io_dram_0_rresp_bits_rdata_14),
    .io_dram_0_rresp_bits_rdata_15(fringeCommon_io_dram_0_rresp_bits_rdata_15),
    .io_dram_0_rresp_bits_tag_streamId(fringeCommon_io_dram_0_rresp_bits_tag_streamId),
    .io_dram_0_wresp_ready(fringeCommon_io_dram_0_wresp_ready),
    .io_dram_0_wresp_valid(fringeCommon_io_dram_0_wresp_valid),
    .io_dram_0_wresp_bits_tag_streamId(fringeCommon_io_dram_0_wresp_bits_tag_streamId),
    .io_dram_1_cmd_ready(fringeCommon_io_dram_1_cmd_ready),
    .io_dram_1_cmd_valid(fringeCommon_io_dram_1_cmd_valid),
    .io_dram_1_cmd_bits_addr(fringeCommon_io_dram_1_cmd_bits_addr),
    .io_dram_1_cmd_bits_size(fringeCommon_io_dram_1_cmd_bits_size),
    .io_dram_1_cmd_bits_isWr(fringeCommon_io_dram_1_cmd_bits_isWr),
    .io_dram_1_cmd_bits_tag_uid(fringeCommon_io_dram_1_cmd_bits_tag_uid),
    .io_dram_1_cmd_bits_tag_streamId(fringeCommon_io_dram_1_cmd_bits_tag_streamId),
    .io_dram_1_wdata_ready(fringeCommon_io_dram_1_wdata_ready),
    .io_dram_1_wdata_valid(fringeCommon_io_dram_1_wdata_valid),
    .io_dram_1_wdata_bits_wdata_0(fringeCommon_io_dram_1_wdata_bits_wdata_0),
    .io_dram_1_wdata_bits_wdata_1(fringeCommon_io_dram_1_wdata_bits_wdata_1),
    .io_dram_1_wdata_bits_wdata_2(fringeCommon_io_dram_1_wdata_bits_wdata_2),
    .io_dram_1_wdata_bits_wdata_3(fringeCommon_io_dram_1_wdata_bits_wdata_3),
    .io_dram_1_wdata_bits_wdata_4(fringeCommon_io_dram_1_wdata_bits_wdata_4),
    .io_dram_1_wdata_bits_wdata_5(fringeCommon_io_dram_1_wdata_bits_wdata_5),
    .io_dram_1_wdata_bits_wdata_6(fringeCommon_io_dram_1_wdata_bits_wdata_6),
    .io_dram_1_wdata_bits_wdata_7(fringeCommon_io_dram_1_wdata_bits_wdata_7),
    .io_dram_1_wdata_bits_wdata_8(fringeCommon_io_dram_1_wdata_bits_wdata_8),
    .io_dram_1_wdata_bits_wdata_9(fringeCommon_io_dram_1_wdata_bits_wdata_9),
    .io_dram_1_wdata_bits_wdata_10(fringeCommon_io_dram_1_wdata_bits_wdata_10),
    .io_dram_1_wdata_bits_wdata_11(fringeCommon_io_dram_1_wdata_bits_wdata_11),
    .io_dram_1_wdata_bits_wdata_12(fringeCommon_io_dram_1_wdata_bits_wdata_12),
    .io_dram_1_wdata_bits_wdata_13(fringeCommon_io_dram_1_wdata_bits_wdata_13),
    .io_dram_1_wdata_bits_wdata_14(fringeCommon_io_dram_1_wdata_bits_wdata_14),
    .io_dram_1_wdata_bits_wdata_15(fringeCommon_io_dram_1_wdata_bits_wdata_15),
    .io_dram_1_wdata_bits_wstrb_0(fringeCommon_io_dram_1_wdata_bits_wstrb_0),
    .io_dram_1_wdata_bits_wstrb_1(fringeCommon_io_dram_1_wdata_bits_wstrb_1),
    .io_dram_1_wdata_bits_wstrb_2(fringeCommon_io_dram_1_wdata_bits_wstrb_2),
    .io_dram_1_wdata_bits_wstrb_3(fringeCommon_io_dram_1_wdata_bits_wstrb_3),
    .io_dram_1_wdata_bits_wstrb_4(fringeCommon_io_dram_1_wdata_bits_wstrb_4),
    .io_dram_1_wdata_bits_wstrb_5(fringeCommon_io_dram_1_wdata_bits_wstrb_5),
    .io_dram_1_wdata_bits_wstrb_6(fringeCommon_io_dram_1_wdata_bits_wstrb_6),
    .io_dram_1_wdata_bits_wstrb_7(fringeCommon_io_dram_1_wdata_bits_wstrb_7),
    .io_dram_1_wdata_bits_wstrb_8(fringeCommon_io_dram_1_wdata_bits_wstrb_8),
    .io_dram_1_wdata_bits_wstrb_9(fringeCommon_io_dram_1_wdata_bits_wstrb_9),
    .io_dram_1_wdata_bits_wstrb_10(fringeCommon_io_dram_1_wdata_bits_wstrb_10),
    .io_dram_1_wdata_bits_wstrb_11(fringeCommon_io_dram_1_wdata_bits_wstrb_11),
    .io_dram_1_wdata_bits_wstrb_12(fringeCommon_io_dram_1_wdata_bits_wstrb_12),
    .io_dram_1_wdata_bits_wstrb_13(fringeCommon_io_dram_1_wdata_bits_wstrb_13),
    .io_dram_1_wdata_bits_wstrb_14(fringeCommon_io_dram_1_wdata_bits_wstrb_14),
    .io_dram_1_wdata_bits_wstrb_15(fringeCommon_io_dram_1_wdata_bits_wstrb_15),
    .io_dram_1_wdata_bits_wstrb_16(fringeCommon_io_dram_1_wdata_bits_wstrb_16),
    .io_dram_1_wdata_bits_wstrb_17(fringeCommon_io_dram_1_wdata_bits_wstrb_17),
    .io_dram_1_wdata_bits_wstrb_18(fringeCommon_io_dram_1_wdata_bits_wstrb_18),
    .io_dram_1_wdata_bits_wstrb_19(fringeCommon_io_dram_1_wdata_bits_wstrb_19),
    .io_dram_1_wdata_bits_wstrb_20(fringeCommon_io_dram_1_wdata_bits_wstrb_20),
    .io_dram_1_wdata_bits_wstrb_21(fringeCommon_io_dram_1_wdata_bits_wstrb_21),
    .io_dram_1_wdata_bits_wstrb_22(fringeCommon_io_dram_1_wdata_bits_wstrb_22),
    .io_dram_1_wdata_bits_wstrb_23(fringeCommon_io_dram_1_wdata_bits_wstrb_23),
    .io_dram_1_wdata_bits_wstrb_24(fringeCommon_io_dram_1_wdata_bits_wstrb_24),
    .io_dram_1_wdata_bits_wstrb_25(fringeCommon_io_dram_1_wdata_bits_wstrb_25),
    .io_dram_1_wdata_bits_wstrb_26(fringeCommon_io_dram_1_wdata_bits_wstrb_26),
    .io_dram_1_wdata_bits_wstrb_27(fringeCommon_io_dram_1_wdata_bits_wstrb_27),
    .io_dram_1_wdata_bits_wstrb_28(fringeCommon_io_dram_1_wdata_bits_wstrb_28),
    .io_dram_1_wdata_bits_wstrb_29(fringeCommon_io_dram_1_wdata_bits_wstrb_29),
    .io_dram_1_wdata_bits_wstrb_30(fringeCommon_io_dram_1_wdata_bits_wstrb_30),
    .io_dram_1_wdata_bits_wstrb_31(fringeCommon_io_dram_1_wdata_bits_wstrb_31),
    .io_dram_1_wdata_bits_wstrb_32(fringeCommon_io_dram_1_wdata_bits_wstrb_32),
    .io_dram_1_wdata_bits_wstrb_33(fringeCommon_io_dram_1_wdata_bits_wstrb_33),
    .io_dram_1_wdata_bits_wstrb_34(fringeCommon_io_dram_1_wdata_bits_wstrb_34),
    .io_dram_1_wdata_bits_wstrb_35(fringeCommon_io_dram_1_wdata_bits_wstrb_35),
    .io_dram_1_wdata_bits_wstrb_36(fringeCommon_io_dram_1_wdata_bits_wstrb_36),
    .io_dram_1_wdata_bits_wstrb_37(fringeCommon_io_dram_1_wdata_bits_wstrb_37),
    .io_dram_1_wdata_bits_wstrb_38(fringeCommon_io_dram_1_wdata_bits_wstrb_38),
    .io_dram_1_wdata_bits_wstrb_39(fringeCommon_io_dram_1_wdata_bits_wstrb_39),
    .io_dram_1_wdata_bits_wstrb_40(fringeCommon_io_dram_1_wdata_bits_wstrb_40),
    .io_dram_1_wdata_bits_wstrb_41(fringeCommon_io_dram_1_wdata_bits_wstrb_41),
    .io_dram_1_wdata_bits_wstrb_42(fringeCommon_io_dram_1_wdata_bits_wstrb_42),
    .io_dram_1_wdata_bits_wstrb_43(fringeCommon_io_dram_1_wdata_bits_wstrb_43),
    .io_dram_1_wdata_bits_wstrb_44(fringeCommon_io_dram_1_wdata_bits_wstrb_44),
    .io_dram_1_wdata_bits_wstrb_45(fringeCommon_io_dram_1_wdata_bits_wstrb_45),
    .io_dram_1_wdata_bits_wstrb_46(fringeCommon_io_dram_1_wdata_bits_wstrb_46),
    .io_dram_1_wdata_bits_wstrb_47(fringeCommon_io_dram_1_wdata_bits_wstrb_47),
    .io_dram_1_wdata_bits_wstrb_48(fringeCommon_io_dram_1_wdata_bits_wstrb_48),
    .io_dram_1_wdata_bits_wstrb_49(fringeCommon_io_dram_1_wdata_bits_wstrb_49),
    .io_dram_1_wdata_bits_wstrb_50(fringeCommon_io_dram_1_wdata_bits_wstrb_50),
    .io_dram_1_wdata_bits_wstrb_51(fringeCommon_io_dram_1_wdata_bits_wstrb_51),
    .io_dram_1_wdata_bits_wstrb_52(fringeCommon_io_dram_1_wdata_bits_wstrb_52),
    .io_dram_1_wdata_bits_wstrb_53(fringeCommon_io_dram_1_wdata_bits_wstrb_53),
    .io_dram_1_wdata_bits_wstrb_54(fringeCommon_io_dram_1_wdata_bits_wstrb_54),
    .io_dram_1_wdata_bits_wstrb_55(fringeCommon_io_dram_1_wdata_bits_wstrb_55),
    .io_dram_1_wdata_bits_wstrb_56(fringeCommon_io_dram_1_wdata_bits_wstrb_56),
    .io_dram_1_wdata_bits_wstrb_57(fringeCommon_io_dram_1_wdata_bits_wstrb_57),
    .io_dram_1_wdata_bits_wstrb_58(fringeCommon_io_dram_1_wdata_bits_wstrb_58),
    .io_dram_1_wdata_bits_wstrb_59(fringeCommon_io_dram_1_wdata_bits_wstrb_59),
    .io_dram_1_wdata_bits_wstrb_60(fringeCommon_io_dram_1_wdata_bits_wstrb_60),
    .io_dram_1_wdata_bits_wstrb_61(fringeCommon_io_dram_1_wdata_bits_wstrb_61),
    .io_dram_1_wdata_bits_wstrb_62(fringeCommon_io_dram_1_wdata_bits_wstrb_62),
    .io_dram_1_wdata_bits_wstrb_63(fringeCommon_io_dram_1_wdata_bits_wstrb_63),
    .io_dram_1_rresp_ready(fringeCommon_io_dram_1_rresp_ready),
    .io_dram_1_rresp_valid(fringeCommon_io_dram_1_rresp_valid),
    .io_dram_1_rresp_bits_rdata_0(fringeCommon_io_dram_1_rresp_bits_rdata_0),
    .io_dram_1_rresp_bits_rdata_1(fringeCommon_io_dram_1_rresp_bits_rdata_1),
    .io_dram_1_rresp_bits_rdata_2(fringeCommon_io_dram_1_rresp_bits_rdata_2),
    .io_dram_1_rresp_bits_rdata_3(fringeCommon_io_dram_1_rresp_bits_rdata_3),
    .io_dram_1_rresp_bits_rdata_4(fringeCommon_io_dram_1_rresp_bits_rdata_4),
    .io_dram_1_rresp_bits_rdata_5(fringeCommon_io_dram_1_rresp_bits_rdata_5),
    .io_dram_1_rresp_bits_rdata_6(fringeCommon_io_dram_1_rresp_bits_rdata_6),
    .io_dram_1_rresp_bits_rdata_7(fringeCommon_io_dram_1_rresp_bits_rdata_7),
    .io_dram_1_rresp_bits_rdata_8(fringeCommon_io_dram_1_rresp_bits_rdata_8),
    .io_dram_1_rresp_bits_rdata_9(fringeCommon_io_dram_1_rresp_bits_rdata_9),
    .io_dram_1_rresp_bits_rdata_10(fringeCommon_io_dram_1_rresp_bits_rdata_10),
    .io_dram_1_rresp_bits_rdata_11(fringeCommon_io_dram_1_rresp_bits_rdata_11),
    .io_dram_1_rresp_bits_rdata_12(fringeCommon_io_dram_1_rresp_bits_rdata_12),
    .io_dram_1_rresp_bits_rdata_13(fringeCommon_io_dram_1_rresp_bits_rdata_13),
    .io_dram_1_rresp_bits_rdata_14(fringeCommon_io_dram_1_rresp_bits_rdata_14),
    .io_dram_1_rresp_bits_rdata_15(fringeCommon_io_dram_1_rresp_bits_rdata_15),
    .io_dram_1_rresp_bits_tag_streamId(fringeCommon_io_dram_1_rresp_bits_tag_streamId),
    .io_dram_1_wresp_ready(fringeCommon_io_dram_1_wresp_ready),
    .io_dram_1_wresp_valid(fringeCommon_io_dram_1_wresp_valid),
    .io_dram_1_wresp_bits_tag_streamId(fringeCommon_io_dram_1_wresp_bits_tag_streamId),
    .io_dram_2_cmd_ready(fringeCommon_io_dram_2_cmd_ready),
    .io_dram_2_cmd_valid(fringeCommon_io_dram_2_cmd_valid),
    .io_dram_2_cmd_bits_addr(fringeCommon_io_dram_2_cmd_bits_addr),
    .io_dram_2_cmd_bits_size(fringeCommon_io_dram_2_cmd_bits_size),
    .io_dram_2_cmd_bits_isWr(fringeCommon_io_dram_2_cmd_bits_isWr),
    .io_dram_2_cmd_bits_tag_uid(fringeCommon_io_dram_2_cmd_bits_tag_uid),
    .io_dram_2_cmd_bits_tag_streamId(fringeCommon_io_dram_2_cmd_bits_tag_streamId),
    .io_dram_2_wdata_ready(fringeCommon_io_dram_2_wdata_ready),
    .io_dram_2_wdata_valid(fringeCommon_io_dram_2_wdata_valid),
    .io_dram_2_wdata_bits_wdata_0(fringeCommon_io_dram_2_wdata_bits_wdata_0),
    .io_dram_2_wdata_bits_wdata_1(fringeCommon_io_dram_2_wdata_bits_wdata_1),
    .io_dram_2_wdata_bits_wdata_2(fringeCommon_io_dram_2_wdata_bits_wdata_2),
    .io_dram_2_wdata_bits_wdata_3(fringeCommon_io_dram_2_wdata_bits_wdata_3),
    .io_dram_2_wdata_bits_wdata_4(fringeCommon_io_dram_2_wdata_bits_wdata_4),
    .io_dram_2_wdata_bits_wdata_5(fringeCommon_io_dram_2_wdata_bits_wdata_5),
    .io_dram_2_wdata_bits_wdata_6(fringeCommon_io_dram_2_wdata_bits_wdata_6),
    .io_dram_2_wdata_bits_wdata_7(fringeCommon_io_dram_2_wdata_bits_wdata_7),
    .io_dram_2_wdata_bits_wdata_8(fringeCommon_io_dram_2_wdata_bits_wdata_8),
    .io_dram_2_wdata_bits_wdata_9(fringeCommon_io_dram_2_wdata_bits_wdata_9),
    .io_dram_2_wdata_bits_wdata_10(fringeCommon_io_dram_2_wdata_bits_wdata_10),
    .io_dram_2_wdata_bits_wdata_11(fringeCommon_io_dram_2_wdata_bits_wdata_11),
    .io_dram_2_wdata_bits_wdata_12(fringeCommon_io_dram_2_wdata_bits_wdata_12),
    .io_dram_2_wdata_bits_wdata_13(fringeCommon_io_dram_2_wdata_bits_wdata_13),
    .io_dram_2_wdata_bits_wdata_14(fringeCommon_io_dram_2_wdata_bits_wdata_14),
    .io_dram_2_wdata_bits_wdata_15(fringeCommon_io_dram_2_wdata_bits_wdata_15),
    .io_dram_2_wdata_bits_wstrb_0(fringeCommon_io_dram_2_wdata_bits_wstrb_0),
    .io_dram_2_wdata_bits_wstrb_1(fringeCommon_io_dram_2_wdata_bits_wstrb_1),
    .io_dram_2_wdata_bits_wstrb_2(fringeCommon_io_dram_2_wdata_bits_wstrb_2),
    .io_dram_2_wdata_bits_wstrb_3(fringeCommon_io_dram_2_wdata_bits_wstrb_3),
    .io_dram_2_wdata_bits_wstrb_4(fringeCommon_io_dram_2_wdata_bits_wstrb_4),
    .io_dram_2_wdata_bits_wstrb_5(fringeCommon_io_dram_2_wdata_bits_wstrb_5),
    .io_dram_2_wdata_bits_wstrb_6(fringeCommon_io_dram_2_wdata_bits_wstrb_6),
    .io_dram_2_wdata_bits_wstrb_7(fringeCommon_io_dram_2_wdata_bits_wstrb_7),
    .io_dram_2_wdata_bits_wstrb_8(fringeCommon_io_dram_2_wdata_bits_wstrb_8),
    .io_dram_2_wdata_bits_wstrb_9(fringeCommon_io_dram_2_wdata_bits_wstrb_9),
    .io_dram_2_wdata_bits_wstrb_10(fringeCommon_io_dram_2_wdata_bits_wstrb_10),
    .io_dram_2_wdata_bits_wstrb_11(fringeCommon_io_dram_2_wdata_bits_wstrb_11),
    .io_dram_2_wdata_bits_wstrb_12(fringeCommon_io_dram_2_wdata_bits_wstrb_12),
    .io_dram_2_wdata_bits_wstrb_13(fringeCommon_io_dram_2_wdata_bits_wstrb_13),
    .io_dram_2_wdata_bits_wstrb_14(fringeCommon_io_dram_2_wdata_bits_wstrb_14),
    .io_dram_2_wdata_bits_wstrb_15(fringeCommon_io_dram_2_wdata_bits_wstrb_15),
    .io_dram_2_wdata_bits_wstrb_16(fringeCommon_io_dram_2_wdata_bits_wstrb_16),
    .io_dram_2_wdata_bits_wstrb_17(fringeCommon_io_dram_2_wdata_bits_wstrb_17),
    .io_dram_2_wdata_bits_wstrb_18(fringeCommon_io_dram_2_wdata_bits_wstrb_18),
    .io_dram_2_wdata_bits_wstrb_19(fringeCommon_io_dram_2_wdata_bits_wstrb_19),
    .io_dram_2_wdata_bits_wstrb_20(fringeCommon_io_dram_2_wdata_bits_wstrb_20),
    .io_dram_2_wdata_bits_wstrb_21(fringeCommon_io_dram_2_wdata_bits_wstrb_21),
    .io_dram_2_wdata_bits_wstrb_22(fringeCommon_io_dram_2_wdata_bits_wstrb_22),
    .io_dram_2_wdata_bits_wstrb_23(fringeCommon_io_dram_2_wdata_bits_wstrb_23),
    .io_dram_2_wdata_bits_wstrb_24(fringeCommon_io_dram_2_wdata_bits_wstrb_24),
    .io_dram_2_wdata_bits_wstrb_25(fringeCommon_io_dram_2_wdata_bits_wstrb_25),
    .io_dram_2_wdata_bits_wstrb_26(fringeCommon_io_dram_2_wdata_bits_wstrb_26),
    .io_dram_2_wdata_bits_wstrb_27(fringeCommon_io_dram_2_wdata_bits_wstrb_27),
    .io_dram_2_wdata_bits_wstrb_28(fringeCommon_io_dram_2_wdata_bits_wstrb_28),
    .io_dram_2_wdata_bits_wstrb_29(fringeCommon_io_dram_2_wdata_bits_wstrb_29),
    .io_dram_2_wdata_bits_wstrb_30(fringeCommon_io_dram_2_wdata_bits_wstrb_30),
    .io_dram_2_wdata_bits_wstrb_31(fringeCommon_io_dram_2_wdata_bits_wstrb_31),
    .io_dram_2_wdata_bits_wstrb_32(fringeCommon_io_dram_2_wdata_bits_wstrb_32),
    .io_dram_2_wdata_bits_wstrb_33(fringeCommon_io_dram_2_wdata_bits_wstrb_33),
    .io_dram_2_wdata_bits_wstrb_34(fringeCommon_io_dram_2_wdata_bits_wstrb_34),
    .io_dram_2_wdata_bits_wstrb_35(fringeCommon_io_dram_2_wdata_bits_wstrb_35),
    .io_dram_2_wdata_bits_wstrb_36(fringeCommon_io_dram_2_wdata_bits_wstrb_36),
    .io_dram_2_wdata_bits_wstrb_37(fringeCommon_io_dram_2_wdata_bits_wstrb_37),
    .io_dram_2_wdata_bits_wstrb_38(fringeCommon_io_dram_2_wdata_bits_wstrb_38),
    .io_dram_2_wdata_bits_wstrb_39(fringeCommon_io_dram_2_wdata_bits_wstrb_39),
    .io_dram_2_wdata_bits_wstrb_40(fringeCommon_io_dram_2_wdata_bits_wstrb_40),
    .io_dram_2_wdata_bits_wstrb_41(fringeCommon_io_dram_2_wdata_bits_wstrb_41),
    .io_dram_2_wdata_bits_wstrb_42(fringeCommon_io_dram_2_wdata_bits_wstrb_42),
    .io_dram_2_wdata_bits_wstrb_43(fringeCommon_io_dram_2_wdata_bits_wstrb_43),
    .io_dram_2_wdata_bits_wstrb_44(fringeCommon_io_dram_2_wdata_bits_wstrb_44),
    .io_dram_2_wdata_bits_wstrb_45(fringeCommon_io_dram_2_wdata_bits_wstrb_45),
    .io_dram_2_wdata_bits_wstrb_46(fringeCommon_io_dram_2_wdata_bits_wstrb_46),
    .io_dram_2_wdata_bits_wstrb_47(fringeCommon_io_dram_2_wdata_bits_wstrb_47),
    .io_dram_2_wdata_bits_wstrb_48(fringeCommon_io_dram_2_wdata_bits_wstrb_48),
    .io_dram_2_wdata_bits_wstrb_49(fringeCommon_io_dram_2_wdata_bits_wstrb_49),
    .io_dram_2_wdata_bits_wstrb_50(fringeCommon_io_dram_2_wdata_bits_wstrb_50),
    .io_dram_2_wdata_bits_wstrb_51(fringeCommon_io_dram_2_wdata_bits_wstrb_51),
    .io_dram_2_wdata_bits_wstrb_52(fringeCommon_io_dram_2_wdata_bits_wstrb_52),
    .io_dram_2_wdata_bits_wstrb_53(fringeCommon_io_dram_2_wdata_bits_wstrb_53),
    .io_dram_2_wdata_bits_wstrb_54(fringeCommon_io_dram_2_wdata_bits_wstrb_54),
    .io_dram_2_wdata_bits_wstrb_55(fringeCommon_io_dram_2_wdata_bits_wstrb_55),
    .io_dram_2_wdata_bits_wstrb_56(fringeCommon_io_dram_2_wdata_bits_wstrb_56),
    .io_dram_2_wdata_bits_wstrb_57(fringeCommon_io_dram_2_wdata_bits_wstrb_57),
    .io_dram_2_wdata_bits_wstrb_58(fringeCommon_io_dram_2_wdata_bits_wstrb_58),
    .io_dram_2_wdata_bits_wstrb_59(fringeCommon_io_dram_2_wdata_bits_wstrb_59),
    .io_dram_2_wdata_bits_wstrb_60(fringeCommon_io_dram_2_wdata_bits_wstrb_60),
    .io_dram_2_wdata_bits_wstrb_61(fringeCommon_io_dram_2_wdata_bits_wstrb_61),
    .io_dram_2_wdata_bits_wstrb_62(fringeCommon_io_dram_2_wdata_bits_wstrb_62),
    .io_dram_2_wdata_bits_wstrb_63(fringeCommon_io_dram_2_wdata_bits_wstrb_63),
    .io_dram_2_rresp_ready(fringeCommon_io_dram_2_rresp_ready),
    .io_dram_2_rresp_valid(fringeCommon_io_dram_2_rresp_valid),
    .io_dram_2_rresp_bits_rdata_0(fringeCommon_io_dram_2_rresp_bits_rdata_0),
    .io_dram_2_rresp_bits_rdata_1(fringeCommon_io_dram_2_rresp_bits_rdata_1),
    .io_dram_2_rresp_bits_rdata_2(fringeCommon_io_dram_2_rresp_bits_rdata_2),
    .io_dram_2_rresp_bits_rdata_3(fringeCommon_io_dram_2_rresp_bits_rdata_3),
    .io_dram_2_rresp_bits_rdata_4(fringeCommon_io_dram_2_rresp_bits_rdata_4),
    .io_dram_2_rresp_bits_rdata_5(fringeCommon_io_dram_2_rresp_bits_rdata_5),
    .io_dram_2_rresp_bits_rdata_6(fringeCommon_io_dram_2_rresp_bits_rdata_6),
    .io_dram_2_rresp_bits_rdata_7(fringeCommon_io_dram_2_rresp_bits_rdata_7),
    .io_dram_2_rresp_bits_rdata_8(fringeCommon_io_dram_2_rresp_bits_rdata_8),
    .io_dram_2_rresp_bits_rdata_9(fringeCommon_io_dram_2_rresp_bits_rdata_9),
    .io_dram_2_rresp_bits_rdata_10(fringeCommon_io_dram_2_rresp_bits_rdata_10),
    .io_dram_2_rresp_bits_rdata_11(fringeCommon_io_dram_2_rresp_bits_rdata_11),
    .io_dram_2_rresp_bits_rdata_12(fringeCommon_io_dram_2_rresp_bits_rdata_12),
    .io_dram_2_rresp_bits_rdata_13(fringeCommon_io_dram_2_rresp_bits_rdata_13),
    .io_dram_2_rresp_bits_rdata_14(fringeCommon_io_dram_2_rresp_bits_rdata_14),
    .io_dram_2_rresp_bits_rdata_15(fringeCommon_io_dram_2_rresp_bits_rdata_15),
    .io_dram_2_rresp_bits_tag_streamId(fringeCommon_io_dram_2_rresp_bits_tag_streamId),
    .io_dram_2_wresp_ready(fringeCommon_io_dram_2_wresp_ready),
    .io_dram_2_wresp_valid(fringeCommon_io_dram_2_wresp_valid),
    .io_dram_2_wresp_bits_tag_streamId(fringeCommon_io_dram_2_wresp_bits_tag_streamId),
    .io_dram_3_cmd_ready(fringeCommon_io_dram_3_cmd_ready),
    .io_dram_3_cmd_valid(fringeCommon_io_dram_3_cmd_valid),
    .io_dram_3_cmd_bits_addr(fringeCommon_io_dram_3_cmd_bits_addr),
    .io_dram_3_cmd_bits_size(fringeCommon_io_dram_3_cmd_bits_size),
    .io_dram_3_cmd_bits_isWr(fringeCommon_io_dram_3_cmd_bits_isWr),
    .io_dram_3_cmd_bits_tag_uid(fringeCommon_io_dram_3_cmd_bits_tag_uid),
    .io_dram_3_cmd_bits_tag_streamId(fringeCommon_io_dram_3_cmd_bits_tag_streamId),
    .io_dram_3_wdata_ready(fringeCommon_io_dram_3_wdata_ready),
    .io_dram_3_wdata_valid(fringeCommon_io_dram_3_wdata_valid),
    .io_dram_3_wdata_bits_wdata_0(fringeCommon_io_dram_3_wdata_bits_wdata_0),
    .io_dram_3_wdata_bits_wdata_1(fringeCommon_io_dram_3_wdata_bits_wdata_1),
    .io_dram_3_wdata_bits_wdata_2(fringeCommon_io_dram_3_wdata_bits_wdata_2),
    .io_dram_3_wdata_bits_wdata_3(fringeCommon_io_dram_3_wdata_bits_wdata_3),
    .io_dram_3_wdata_bits_wdata_4(fringeCommon_io_dram_3_wdata_bits_wdata_4),
    .io_dram_3_wdata_bits_wdata_5(fringeCommon_io_dram_3_wdata_bits_wdata_5),
    .io_dram_3_wdata_bits_wdata_6(fringeCommon_io_dram_3_wdata_bits_wdata_6),
    .io_dram_3_wdata_bits_wdata_7(fringeCommon_io_dram_3_wdata_bits_wdata_7),
    .io_dram_3_wdata_bits_wdata_8(fringeCommon_io_dram_3_wdata_bits_wdata_8),
    .io_dram_3_wdata_bits_wdata_9(fringeCommon_io_dram_3_wdata_bits_wdata_9),
    .io_dram_3_wdata_bits_wdata_10(fringeCommon_io_dram_3_wdata_bits_wdata_10),
    .io_dram_3_wdata_bits_wdata_11(fringeCommon_io_dram_3_wdata_bits_wdata_11),
    .io_dram_3_wdata_bits_wdata_12(fringeCommon_io_dram_3_wdata_bits_wdata_12),
    .io_dram_3_wdata_bits_wdata_13(fringeCommon_io_dram_3_wdata_bits_wdata_13),
    .io_dram_3_wdata_bits_wdata_14(fringeCommon_io_dram_3_wdata_bits_wdata_14),
    .io_dram_3_wdata_bits_wdata_15(fringeCommon_io_dram_3_wdata_bits_wdata_15),
    .io_dram_3_wdata_bits_wstrb_0(fringeCommon_io_dram_3_wdata_bits_wstrb_0),
    .io_dram_3_wdata_bits_wstrb_1(fringeCommon_io_dram_3_wdata_bits_wstrb_1),
    .io_dram_3_wdata_bits_wstrb_2(fringeCommon_io_dram_3_wdata_bits_wstrb_2),
    .io_dram_3_wdata_bits_wstrb_3(fringeCommon_io_dram_3_wdata_bits_wstrb_3),
    .io_dram_3_wdata_bits_wstrb_4(fringeCommon_io_dram_3_wdata_bits_wstrb_4),
    .io_dram_3_wdata_bits_wstrb_5(fringeCommon_io_dram_3_wdata_bits_wstrb_5),
    .io_dram_3_wdata_bits_wstrb_6(fringeCommon_io_dram_3_wdata_bits_wstrb_6),
    .io_dram_3_wdata_bits_wstrb_7(fringeCommon_io_dram_3_wdata_bits_wstrb_7),
    .io_dram_3_wdata_bits_wstrb_8(fringeCommon_io_dram_3_wdata_bits_wstrb_8),
    .io_dram_3_wdata_bits_wstrb_9(fringeCommon_io_dram_3_wdata_bits_wstrb_9),
    .io_dram_3_wdata_bits_wstrb_10(fringeCommon_io_dram_3_wdata_bits_wstrb_10),
    .io_dram_3_wdata_bits_wstrb_11(fringeCommon_io_dram_3_wdata_bits_wstrb_11),
    .io_dram_3_wdata_bits_wstrb_12(fringeCommon_io_dram_3_wdata_bits_wstrb_12),
    .io_dram_3_wdata_bits_wstrb_13(fringeCommon_io_dram_3_wdata_bits_wstrb_13),
    .io_dram_3_wdata_bits_wstrb_14(fringeCommon_io_dram_3_wdata_bits_wstrb_14),
    .io_dram_3_wdata_bits_wstrb_15(fringeCommon_io_dram_3_wdata_bits_wstrb_15),
    .io_dram_3_wdata_bits_wstrb_16(fringeCommon_io_dram_3_wdata_bits_wstrb_16),
    .io_dram_3_wdata_bits_wstrb_17(fringeCommon_io_dram_3_wdata_bits_wstrb_17),
    .io_dram_3_wdata_bits_wstrb_18(fringeCommon_io_dram_3_wdata_bits_wstrb_18),
    .io_dram_3_wdata_bits_wstrb_19(fringeCommon_io_dram_3_wdata_bits_wstrb_19),
    .io_dram_3_wdata_bits_wstrb_20(fringeCommon_io_dram_3_wdata_bits_wstrb_20),
    .io_dram_3_wdata_bits_wstrb_21(fringeCommon_io_dram_3_wdata_bits_wstrb_21),
    .io_dram_3_wdata_bits_wstrb_22(fringeCommon_io_dram_3_wdata_bits_wstrb_22),
    .io_dram_3_wdata_bits_wstrb_23(fringeCommon_io_dram_3_wdata_bits_wstrb_23),
    .io_dram_3_wdata_bits_wstrb_24(fringeCommon_io_dram_3_wdata_bits_wstrb_24),
    .io_dram_3_wdata_bits_wstrb_25(fringeCommon_io_dram_3_wdata_bits_wstrb_25),
    .io_dram_3_wdata_bits_wstrb_26(fringeCommon_io_dram_3_wdata_bits_wstrb_26),
    .io_dram_3_wdata_bits_wstrb_27(fringeCommon_io_dram_3_wdata_bits_wstrb_27),
    .io_dram_3_wdata_bits_wstrb_28(fringeCommon_io_dram_3_wdata_bits_wstrb_28),
    .io_dram_3_wdata_bits_wstrb_29(fringeCommon_io_dram_3_wdata_bits_wstrb_29),
    .io_dram_3_wdata_bits_wstrb_30(fringeCommon_io_dram_3_wdata_bits_wstrb_30),
    .io_dram_3_wdata_bits_wstrb_31(fringeCommon_io_dram_3_wdata_bits_wstrb_31),
    .io_dram_3_wdata_bits_wstrb_32(fringeCommon_io_dram_3_wdata_bits_wstrb_32),
    .io_dram_3_wdata_bits_wstrb_33(fringeCommon_io_dram_3_wdata_bits_wstrb_33),
    .io_dram_3_wdata_bits_wstrb_34(fringeCommon_io_dram_3_wdata_bits_wstrb_34),
    .io_dram_3_wdata_bits_wstrb_35(fringeCommon_io_dram_3_wdata_bits_wstrb_35),
    .io_dram_3_wdata_bits_wstrb_36(fringeCommon_io_dram_3_wdata_bits_wstrb_36),
    .io_dram_3_wdata_bits_wstrb_37(fringeCommon_io_dram_3_wdata_bits_wstrb_37),
    .io_dram_3_wdata_bits_wstrb_38(fringeCommon_io_dram_3_wdata_bits_wstrb_38),
    .io_dram_3_wdata_bits_wstrb_39(fringeCommon_io_dram_3_wdata_bits_wstrb_39),
    .io_dram_3_wdata_bits_wstrb_40(fringeCommon_io_dram_3_wdata_bits_wstrb_40),
    .io_dram_3_wdata_bits_wstrb_41(fringeCommon_io_dram_3_wdata_bits_wstrb_41),
    .io_dram_3_wdata_bits_wstrb_42(fringeCommon_io_dram_3_wdata_bits_wstrb_42),
    .io_dram_3_wdata_bits_wstrb_43(fringeCommon_io_dram_3_wdata_bits_wstrb_43),
    .io_dram_3_wdata_bits_wstrb_44(fringeCommon_io_dram_3_wdata_bits_wstrb_44),
    .io_dram_3_wdata_bits_wstrb_45(fringeCommon_io_dram_3_wdata_bits_wstrb_45),
    .io_dram_3_wdata_bits_wstrb_46(fringeCommon_io_dram_3_wdata_bits_wstrb_46),
    .io_dram_3_wdata_bits_wstrb_47(fringeCommon_io_dram_3_wdata_bits_wstrb_47),
    .io_dram_3_wdata_bits_wstrb_48(fringeCommon_io_dram_3_wdata_bits_wstrb_48),
    .io_dram_3_wdata_bits_wstrb_49(fringeCommon_io_dram_3_wdata_bits_wstrb_49),
    .io_dram_3_wdata_bits_wstrb_50(fringeCommon_io_dram_3_wdata_bits_wstrb_50),
    .io_dram_3_wdata_bits_wstrb_51(fringeCommon_io_dram_3_wdata_bits_wstrb_51),
    .io_dram_3_wdata_bits_wstrb_52(fringeCommon_io_dram_3_wdata_bits_wstrb_52),
    .io_dram_3_wdata_bits_wstrb_53(fringeCommon_io_dram_3_wdata_bits_wstrb_53),
    .io_dram_3_wdata_bits_wstrb_54(fringeCommon_io_dram_3_wdata_bits_wstrb_54),
    .io_dram_3_wdata_bits_wstrb_55(fringeCommon_io_dram_3_wdata_bits_wstrb_55),
    .io_dram_3_wdata_bits_wstrb_56(fringeCommon_io_dram_3_wdata_bits_wstrb_56),
    .io_dram_3_wdata_bits_wstrb_57(fringeCommon_io_dram_3_wdata_bits_wstrb_57),
    .io_dram_3_wdata_bits_wstrb_58(fringeCommon_io_dram_3_wdata_bits_wstrb_58),
    .io_dram_3_wdata_bits_wstrb_59(fringeCommon_io_dram_3_wdata_bits_wstrb_59),
    .io_dram_3_wdata_bits_wstrb_60(fringeCommon_io_dram_3_wdata_bits_wstrb_60),
    .io_dram_3_wdata_bits_wstrb_61(fringeCommon_io_dram_3_wdata_bits_wstrb_61),
    .io_dram_3_wdata_bits_wstrb_62(fringeCommon_io_dram_3_wdata_bits_wstrb_62),
    .io_dram_3_wdata_bits_wstrb_63(fringeCommon_io_dram_3_wdata_bits_wstrb_63),
    .io_dram_3_rresp_ready(fringeCommon_io_dram_3_rresp_ready),
    .io_dram_3_rresp_valid(fringeCommon_io_dram_3_rresp_valid),
    .io_dram_3_rresp_bits_rdata_0(fringeCommon_io_dram_3_rresp_bits_rdata_0),
    .io_dram_3_rresp_bits_rdata_1(fringeCommon_io_dram_3_rresp_bits_rdata_1),
    .io_dram_3_rresp_bits_rdata_2(fringeCommon_io_dram_3_rresp_bits_rdata_2),
    .io_dram_3_rresp_bits_rdata_3(fringeCommon_io_dram_3_rresp_bits_rdata_3),
    .io_dram_3_rresp_bits_rdata_4(fringeCommon_io_dram_3_rresp_bits_rdata_4),
    .io_dram_3_rresp_bits_rdata_5(fringeCommon_io_dram_3_rresp_bits_rdata_5),
    .io_dram_3_rresp_bits_rdata_6(fringeCommon_io_dram_3_rresp_bits_rdata_6),
    .io_dram_3_rresp_bits_rdata_7(fringeCommon_io_dram_3_rresp_bits_rdata_7),
    .io_dram_3_rresp_bits_rdata_8(fringeCommon_io_dram_3_rresp_bits_rdata_8),
    .io_dram_3_rresp_bits_rdata_9(fringeCommon_io_dram_3_rresp_bits_rdata_9),
    .io_dram_3_rresp_bits_rdata_10(fringeCommon_io_dram_3_rresp_bits_rdata_10),
    .io_dram_3_rresp_bits_rdata_11(fringeCommon_io_dram_3_rresp_bits_rdata_11),
    .io_dram_3_rresp_bits_rdata_12(fringeCommon_io_dram_3_rresp_bits_rdata_12),
    .io_dram_3_rresp_bits_rdata_13(fringeCommon_io_dram_3_rresp_bits_rdata_13),
    .io_dram_3_rresp_bits_rdata_14(fringeCommon_io_dram_3_rresp_bits_rdata_14),
    .io_dram_3_rresp_bits_rdata_15(fringeCommon_io_dram_3_rresp_bits_rdata_15),
    .io_dram_3_rresp_bits_tag_streamId(fringeCommon_io_dram_3_rresp_bits_tag_streamId),
    .io_dram_3_wresp_ready(fringeCommon_io_dram_3_wresp_ready),
    .io_dram_3_wresp_valid(fringeCommon_io_dram_3_wresp_valid),
    .io_dram_3_wresp_bits_tag_streamId(fringeCommon_io_dram_3_wresp_bits_tag_streamId),
    .io_TOP_AXI_AWADDR(fringeCommon_io_TOP_AXI_AWADDR),
    .io_TOP_AXI_AWLEN(fringeCommon_io_TOP_AXI_AWLEN),
    .io_TOP_AXI_AWVALID(fringeCommon_io_TOP_AXI_AWVALID),
    .io_TOP_AXI_AWREADY(fringeCommon_io_TOP_AXI_AWREADY),
    .io_TOP_AXI_ARID(fringeCommon_io_TOP_AXI_ARID),
    .io_TOP_AXI_ARADDR(fringeCommon_io_TOP_AXI_ARADDR),
    .io_TOP_AXI_ARLEN(fringeCommon_io_TOP_AXI_ARLEN),
    .io_TOP_AXI_ARSIZE(fringeCommon_io_TOP_AXI_ARSIZE),
    .io_TOP_AXI_ARBURST(fringeCommon_io_TOP_AXI_ARBURST),
    .io_TOP_AXI_ARVALID(fringeCommon_io_TOP_AXI_ARVALID),
    .io_TOP_AXI_ARREADY(fringeCommon_io_TOP_AXI_ARREADY),
    .io_TOP_AXI_WDATA(fringeCommon_io_TOP_AXI_WDATA),
    .io_TOP_AXI_WSTRB(fringeCommon_io_TOP_AXI_WSTRB),
    .io_TOP_AXI_WVALID(fringeCommon_io_TOP_AXI_WVALID),
    .io_TOP_AXI_WREADY(fringeCommon_io_TOP_AXI_WREADY),
    .io_TOP_AXI_RVALID(fringeCommon_io_TOP_AXI_RVALID),
    .io_TOP_AXI_RREADY(fringeCommon_io_TOP_AXI_RREADY),
    .io_TOP_AXI_BVALID(fringeCommon_io_TOP_AXI_BVALID),
    .io_TOP_AXI_BREADY(fringeCommon_io_TOP_AXI_BREADY),
    .io_DWIDTH_AXI_AWADDR(fringeCommon_io_DWIDTH_AXI_AWADDR),
    .io_DWIDTH_AXI_AWLEN(fringeCommon_io_DWIDTH_AXI_AWLEN),
    .io_DWIDTH_AXI_AWVALID(fringeCommon_io_DWIDTH_AXI_AWVALID),
    .io_DWIDTH_AXI_AWREADY(fringeCommon_io_DWIDTH_AXI_AWREADY),
    .io_DWIDTH_AXI_ARADDR(fringeCommon_io_DWIDTH_AXI_ARADDR),
    .io_DWIDTH_AXI_ARLEN(fringeCommon_io_DWIDTH_AXI_ARLEN),
    .io_DWIDTH_AXI_ARSIZE(fringeCommon_io_DWIDTH_AXI_ARSIZE),
    .io_DWIDTH_AXI_ARBURST(fringeCommon_io_DWIDTH_AXI_ARBURST),
    .io_DWIDTH_AXI_ARVALID(fringeCommon_io_DWIDTH_AXI_ARVALID),
    .io_DWIDTH_AXI_ARREADY(fringeCommon_io_DWIDTH_AXI_ARREADY),
    .io_DWIDTH_AXI_WDATA(fringeCommon_io_DWIDTH_AXI_WDATA),
    .io_DWIDTH_AXI_WSTRB(fringeCommon_io_DWIDTH_AXI_WSTRB),
    .io_DWIDTH_AXI_WVALID(fringeCommon_io_DWIDTH_AXI_WVALID),
    .io_DWIDTH_AXI_WREADY(fringeCommon_io_DWIDTH_AXI_WREADY),
    .io_DWIDTH_AXI_RVALID(fringeCommon_io_DWIDTH_AXI_RVALID),
    .io_DWIDTH_AXI_RREADY(fringeCommon_io_DWIDTH_AXI_RREADY),
    .io_DWIDTH_AXI_BVALID(fringeCommon_io_DWIDTH_AXI_BVALID),
    .io_DWIDTH_AXI_BREADY(fringeCommon_io_DWIDTH_AXI_BREADY)
  );
  AXI4LiteToRFBridge AXI4LiteToRFBridge (
    .clock(AXI4LiteToRFBridge_clock),
    .reset(AXI4LiteToRFBridge_reset),
    .io_S_AXI_AWADDR(AXI4LiteToRFBridge_io_S_AXI_AWADDR),
    .io_S_AXI_AWPROT(AXI4LiteToRFBridge_io_S_AXI_AWPROT),
    .io_S_AXI_AWVALID(AXI4LiteToRFBridge_io_S_AXI_AWVALID),
    .io_S_AXI_AWREADY(AXI4LiteToRFBridge_io_S_AXI_AWREADY),
    .io_S_AXI_ARADDR(AXI4LiteToRFBridge_io_S_AXI_ARADDR),
    .io_S_AXI_ARPROT(AXI4LiteToRFBridge_io_S_AXI_ARPROT),
    .io_S_AXI_ARVALID(AXI4LiteToRFBridge_io_S_AXI_ARVALID),
    .io_S_AXI_ARREADY(AXI4LiteToRFBridge_io_S_AXI_ARREADY),
    .io_S_AXI_WDATA(AXI4LiteToRFBridge_io_S_AXI_WDATA),
    .io_S_AXI_WSTRB(AXI4LiteToRFBridge_io_S_AXI_WSTRB),
    .io_S_AXI_WVALID(AXI4LiteToRFBridge_io_S_AXI_WVALID),
    .io_S_AXI_WREADY(AXI4LiteToRFBridge_io_S_AXI_WREADY),
    .io_S_AXI_RDATA(AXI4LiteToRFBridge_io_S_AXI_RDATA),
    .io_S_AXI_RRESP(AXI4LiteToRFBridge_io_S_AXI_RRESP),
    .io_S_AXI_RVALID(AXI4LiteToRFBridge_io_S_AXI_RVALID),
    .io_S_AXI_RREADY(AXI4LiteToRFBridge_io_S_AXI_RREADY),
    .io_S_AXI_BRESP(AXI4LiteToRFBridge_io_S_AXI_BRESP),
    .io_S_AXI_BVALID(AXI4LiteToRFBridge_io_S_AXI_BVALID),
    .io_S_AXI_BREADY(AXI4LiteToRFBridge_io_S_AXI_BREADY),
    .io_raddr(AXI4LiteToRFBridge_io_raddr),
    .io_wen(AXI4LiteToRFBridge_io_wen),
    .io_waddr(AXI4LiteToRFBridge_io_waddr),
    .io_wdata(AXI4LiteToRFBridge_io_wdata),
    .io_rdata(AXI4LiteToRFBridge_io_rdata)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge (
    .io_in_cmd_ready(MAGToAXI4Bridge_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag_uid(MAGToAXI4Bridge_io_in_cmd_bits_tag_uid),
    .io_in_cmd_bits_tag_streamId(MAGToAXI4Bridge_io_in_cmd_bits_tag_streamId),
    .io_in_wdata_ready(MAGToAXI4Bridge_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(MAGToAXI4Bridge_io_in_rresp_ready),
    .io_in_rresp_valid(MAGToAXI4Bridge_io_in_rresp_valid),
    .io_in_rresp_bits_rdata_0(MAGToAXI4Bridge_io_in_rresp_bits_rdata_0),
    .io_in_rresp_bits_rdata_1(MAGToAXI4Bridge_io_in_rresp_bits_rdata_1),
    .io_in_rresp_bits_rdata_2(MAGToAXI4Bridge_io_in_rresp_bits_rdata_2),
    .io_in_rresp_bits_rdata_3(MAGToAXI4Bridge_io_in_rresp_bits_rdata_3),
    .io_in_rresp_bits_rdata_4(MAGToAXI4Bridge_io_in_rresp_bits_rdata_4),
    .io_in_rresp_bits_rdata_5(MAGToAXI4Bridge_io_in_rresp_bits_rdata_5),
    .io_in_rresp_bits_rdata_6(MAGToAXI4Bridge_io_in_rresp_bits_rdata_6),
    .io_in_rresp_bits_rdata_7(MAGToAXI4Bridge_io_in_rresp_bits_rdata_7),
    .io_in_rresp_bits_rdata_8(MAGToAXI4Bridge_io_in_rresp_bits_rdata_8),
    .io_in_rresp_bits_rdata_9(MAGToAXI4Bridge_io_in_rresp_bits_rdata_9),
    .io_in_rresp_bits_rdata_10(MAGToAXI4Bridge_io_in_rresp_bits_rdata_10),
    .io_in_rresp_bits_rdata_11(MAGToAXI4Bridge_io_in_rresp_bits_rdata_11),
    .io_in_rresp_bits_rdata_12(MAGToAXI4Bridge_io_in_rresp_bits_rdata_12),
    .io_in_rresp_bits_rdata_13(MAGToAXI4Bridge_io_in_rresp_bits_rdata_13),
    .io_in_rresp_bits_rdata_14(MAGToAXI4Bridge_io_in_rresp_bits_rdata_14),
    .io_in_rresp_bits_rdata_15(MAGToAXI4Bridge_io_in_rresp_bits_rdata_15),
    .io_in_rresp_bits_tag_streamId(MAGToAXI4Bridge_io_in_rresp_bits_tag_streamId),
    .io_in_wresp_ready(MAGToAXI4Bridge_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_io_in_wresp_valid),
    .io_in_wresp_bits_tag_streamId(MAGToAXI4Bridge_io_in_wresp_bits_tag_streamId),
    .io_M_AXI_AWID(MAGToAXI4Bridge_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_io_M_AXI_WSTRB),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_io_M_AXI_WREADY),
    .io_M_AXI_RID(MAGToAXI4Bridge_io_M_AXI_RID),
    .io_M_AXI_RDATA(MAGToAXI4Bridge_io_M_AXI_RDATA),
    .io_M_AXI_RVALID(MAGToAXI4Bridge_io_M_AXI_RVALID),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_io_M_AXI_BREADY)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge_1 (
    .io_in_cmd_ready(MAGToAXI4Bridge_1_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_1_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_1_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_1_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_1_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag_uid(MAGToAXI4Bridge_1_io_in_cmd_bits_tag_uid),
    .io_in_cmd_bits_tag_streamId(MAGToAXI4Bridge_1_io_in_cmd_bits_tag_streamId),
    .io_in_wdata_ready(MAGToAXI4Bridge_1_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_1_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(MAGToAXI4Bridge_1_io_in_rresp_ready),
    .io_in_rresp_valid(MAGToAXI4Bridge_1_io_in_rresp_valid),
    .io_in_rresp_bits_rdata_0(MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_0),
    .io_in_rresp_bits_rdata_1(MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_1),
    .io_in_rresp_bits_rdata_2(MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_2),
    .io_in_rresp_bits_rdata_3(MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_3),
    .io_in_rresp_bits_rdata_4(MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_4),
    .io_in_rresp_bits_rdata_5(MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_5),
    .io_in_rresp_bits_rdata_6(MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_6),
    .io_in_rresp_bits_rdata_7(MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_7),
    .io_in_rresp_bits_rdata_8(MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_8),
    .io_in_rresp_bits_rdata_9(MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_9),
    .io_in_rresp_bits_rdata_10(MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_10),
    .io_in_rresp_bits_rdata_11(MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_11),
    .io_in_rresp_bits_rdata_12(MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_12),
    .io_in_rresp_bits_rdata_13(MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_13),
    .io_in_rresp_bits_rdata_14(MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_14),
    .io_in_rresp_bits_rdata_15(MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_15),
    .io_in_rresp_bits_tag_streamId(MAGToAXI4Bridge_1_io_in_rresp_bits_tag_streamId),
    .io_in_wresp_ready(MAGToAXI4Bridge_1_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_1_io_in_wresp_valid),
    .io_in_wresp_bits_tag_streamId(MAGToAXI4Bridge_1_io_in_wresp_bits_tag_streamId),
    .io_M_AXI_AWID(MAGToAXI4Bridge_1_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_1_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_1_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_1_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_1_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_1_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_1_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_1_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_1_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_1_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_1_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_1_io_M_AXI_WSTRB),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_1_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_1_io_M_AXI_WREADY),
    .io_M_AXI_RID(MAGToAXI4Bridge_1_io_M_AXI_RID),
    .io_M_AXI_RDATA(MAGToAXI4Bridge_1_io_M_AXI_RDATA),
    .io_M_AXI_RVALID(MAGToAXI4Bridge_1_io_M_AXI_RVALID),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_1_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_1_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_1_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_1_io_M_AXI_BREADY)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge_2 (
    .io_in_cmd_ready(MAGToAXI4Bridge_2_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_2_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_2_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_2_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_2_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag_uid(MAGToAXI4Bridge_2_io_in_cmd_bits_tag_uid),
    .io_in_cmd_bits_tag_streamId(MAGToAXI4Bridge_2_io_in_cmd_bits_tag_streamId),
    .io_in_wdata_ready(MAGToAXI4Bridge_2_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_2_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(MAGToAXI4Bridge_2_io_in_rresp_ready),
    .io_in_rresp_valid(MAGToAXI4Bridge_2_io_in_rresp_valid),
    .io_in_rresp_bits_rdata_0(MAGToAXI4Bridge_2_io_in_rresp_bits_rdata_0),
    .io_in_rresp_bits_rdata_1(MAGToAXI4Bridge_2_io_in_rresp_bits_rdata_1),
    .io_in_rresp_bits_rdata_2(MAGToAXI4Bridge_2_io_in_rresp_bits_rdata_2),
    .io_in_rresp_bits_rdata_3(MAGToAXI4Bridge_2_io_in_rresp_bits_rdata_3),
    .io_in_rresp_bits_rdata_4(MAGToAXI4Bridge_2_io_in_rresp_bits_rdata_4),
    .io_in_rresp_bits_rdata_5(MAGToAXI4Bridge_2_io_in_rresp_bits_rdata_5),
    .io_in_rresp_bits_rdata_6(MAGToAXI4Bridge_2_io_in_rresp_bits_rdata_6),
    .io_in_rresp_bits_rdata_7(MAGToAXI4Bridge_2_io_in_rresp_bits_rdata_7),
    .io_in_rresp_bits_rdata_8(MAGToAXI4Bridge_2_io_in_rresp_bits_rdata_8),
    .io_in_rresp_bits_rdata_9(MAGToAXI4Bridge_2_io_in_rresp_bits_rdata_9),
    .io_in_rresp_bits_rdata_10(MAGToAXI4Bridge_2_io_in_rresp_bits_rdata_10),
    .io_in_rresp_bits_rdata_11(MAGToAXI4Bridge_2_io_in_rresp_bits_rdata_11),
    .io_in_rresp_bits_rdata_12(MAGToAXI4Bridge_2_io_in_rresp_bits_rdata_12),
    .io_in_rresp_bits_rdata_13(MAGToAXI4Bridge_2_io_in_rresp_bits_rdata_13),
    .io_in_rresp_bits_rdata_14(MAGToAXI4Bridge_2_io_in_rresp_bits_rdata_14),
    .io_in_rresp_bits_rdata_15(MAGToAXI4Bridge_2_io_in_rresp_bits_rdata_15),
    .io_in_rresp_bits_tag_streamId(MAGToAXI4Bridge_2_io_in_rresp_bits_tag_streamId),
    .io_in_wresp_ready(MAGToAXI4Bridge_2_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_2_io_in_wresp_valid),
    .io_in_wresp_bits_tag_streamId(MAGToAXI4Bridge_2_io_in_wresp_bits_tag_streamId),
    .io_M_AXI_AWID(MAGToAXI4Bridge_2_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_2_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_2_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_2_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_2_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_2_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_2_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_2_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_2_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_2_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_2_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_2_io_M_AXI_WSTRB),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_2_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_2_io_M_AXI_WREADY),
    .io_M_AXI_RID(MAGToAXI4Bridge_2_io_M_AXI_RID),
    .io_M_AXI_RDATA(MAGToAXI4Bridge_2_io_M_AXI_RDATA),
    .io_M_AXI_RVALID(MAGToAXI4Bridge_2_io_M_AXI_RVALID),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_2_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_2_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_2_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_2_io_M_AXI_BREADY)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge_3 (
    .io_in_cmd_ready(MAGToAXI4Bridge_3_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_3_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_3_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_3_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_3_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag_uid(MAGToAXI4Bridge_3_io_in_cmd_bits_tag_uid),
    .io_in_cmd_bits_tag_streamId(MAGToAXI4Bridge_3_io_in_cmd_bits_tag_streamId),
    .io_in_wdata_ready(MAGToAXI4Bridge_3_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_3_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(MAGToAXI4Bridge_3_io_in_rresp_ready),
    .io_in_rresp_valid(MAGToAXI4Bridge_3_io_in_rresp_valid),
    .io_in_rresp_bits_rdata_0(MAGToAXI4Bridge_3_io_in_rresp_bits_rdata_0),
    .io_in_rresp_bits_rdata_1(MAGToAXI4Bridge_3_io_in_rresp_bits_rdata_1),
    .io_in_rresp_bits_rdata_2(MAGToAXI4Bridge_3_io_in_rresp_bits_rdata_2),
    .io_in_rresp_bits_rdata_3(MAGToAXI4Bridge_3_io_in_rresp_bits_rdata_3),
    .io_in_rresp_bits_rdata_4(MAGToAXI4Bridge_3_io_in_rresp_bits_rdata_4),
    .io_in_rresp_bits_rdata_5(MAGToAXI4Bridge_3_io_in_rresp_bits_rdata_5),
    .io_in_rresp_bits_rdata_6(MAGToAXI4Bridge_3_io_in_rresp_bits_rdata_6),
    .io_in_rresp_bits_rdata_7(MAGToAXI4Bridge_3_io_in_rresp_bits_rdata_7),
    .io_in_rresp_bits_rdata_8(MAGToAXI4Bridge_3_io_in_rresp_bits_rdata_8),
    .io_in_rresp_bits_rdata_9(MAGToAXI4Bridge_3_io_in_rresp_bits_rdata_9),
    .io_in_rresp_bits_rdata_10(MAGToAXI4Bridge_3_io_in_rresp_bits_rdata_10),
    .io_in_rresp_bits_rdata_11(MAGToAXI4Bridge_3_io_in_rresp_bits_rdata_11),
    .io_in_rresp_bits_rdata_12(MAGToAXI4Bridge_3_io_in_rresp_bits_rdata_12),
    .io_in_rresp_bits_rdata_13(MAGToAXI4Bridge_3_io_in_rresp_bits_rdata_13),
    .io_in_rresp_bits_rdata_14(MAGToAXI4Bridge_3_io_in_rresp_bits_rdata_14),
    .io_in_rresp_bits_rdata_15(MAGToAXI4Bridge_3_io_in_rresp_bits_rdata_15),
    .io_in_rresp_bits_tag_streamId(MAGToAXI4Bridge_3_io_in_rresp_bits_tag_streamId),
    .io_in_wresp_ready(MAGToAXI4Bridge_3_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_3_io_in_wresp_valid),
    .io_in_wresp_bits_tag_streamId(MAGToAXI4Bridge_3_io_in_wresp_bits_tag_streamId),
    .io_M_AXI_AWID(MAGToAXI4Bridge_3_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_3_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_3_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_3_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_3_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_3_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_3_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_3_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_3_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_3_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_3_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_3_io_M_AXI_WSTRB),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_3_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_3_io_M_AXI_WREADY),
    .io_M_AXI_RID(MAGToAXI4Bridge_3_io_M_AXI_RID),
    .io_M_AXI_RDATA(MAGToAXI4Bridge_3_io_M_AXI_RDATA),
    .io_M_AXI_RVALID(MAGToAXI4Bridge_3_io_M_AXI_RVALID),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_3_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_3_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_3_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_3_io_M_AXI_BREADY)
  );
  assign io_S_AXI_AWREADY = AXI4LiteToRFBridge_io_S_AXI_AWREADY;
  assign io_S_AXI_ARREADY = AXI4LiteToRFBridge_io_S_AXI_ARREADY;
  assign io_S_AXI_WREADY = AXI4LiteToRFBridge_io_S_AXI_WREADY;
  assign io_S_AXI_RDATA = AXI4LiteToRFBridge_io_S_AXI_RDATA;
  assign io_S_AXI_RRESP = AXI4LiteToRFBridge_io_S_AXI_RRESP;
  assign io_S_AXI_RVALID = AXI4LiteToRFBridge_io_S_AXI_RVALID;
  assign io_S_AXI_BRESP = AXI4LiteToRFBridge_io_S_AXI_BRESP;
  assign io_S_AXI_BVALID = AXI4LiteToRFBridge_io_S_AXI_BVALID;
  assign io_M_AXI_0_AWID = MAGToAXI4Bridge_io_M_AXI_AWID;
  assign io_M_AXI_0_AWADDR = MAGToAXI4Bridge_io_M_AXI_AWADDR;
  assign io_M_AXI_0_AWLEN = MAGToAXI4Bridge_io_M_AXI_AWLEN;
  assign io_M_AXI_0_AWVALID = MAGToAXI4Bridge_io_M_AXI_AWVALID;
  assign io_M_AXI_0_ARID = MAGToAXI4Bridge_io_M_AXI_ARID;
  assign io_M_AXI_0_ARADDR = MAGToAXI4Bridge_io_M_AXI_ARADDR;
  assign io_M_AXI_0_ARLEN = MAGToAXI4Bridge_io_M_AXI_ARLEN;
  assign io_M_AXI_0_ARVALID = MAGToAXI4Bridge_io_M_AXI_ARVALID;
  assign io_M_AXI_0_WDATA = MAGToAXI4Bridge_io_M_AXI_WDATA;
  assign io_M_AXI_0_WSTRB = MAGToAXI4Bridge_io_M_AXI_WSTRB;
  assign io_M_AXI_0_WVALID = MAGToAXI4Bridge_io_M_AXI_WVALID;
  assign io_M_AXI_0_RREADY = MAGToAXI4Bridge_io_M_AXI_RREADY;
  assign io_M_AXI_0_BREADY = MAGToAXI4Bridge_io_M_AXI_BREADY;
  assign io_M_AXI_1_AWID = MAGToAXI4Bridge_1_io_M_AXI_AWID;
  assign io_M_AXI_1_AWADDR = MAGToAXI4Bridge_1_io_M_AXI_AWADDR;
  assign io_M_AXI_1_AWLEN = MAGToAXI4Bridge_1_io_M_AXI_AWLEN;
  assign io_M_AXI_1_AWVALID = MAGToAXI4Bridge_1_io_M_AXI_AWVALID;
  assign io_M_AXI_1_ARID = MAGToAXI4Bridge_1_io_M_AXI_ARID;
  assign io_M_AXI_1_ARADDR = MAGToAXI4Bridge_1_io_M_AXI_ARADDR;
  assign io_M_AXI_1_ARLEN = MAGToAXI4Bridge_1_io_M_AXI_ARLEN;
  assign io_M_AXI_1_ARVALID = MAGToAXI4Bridge_1_io_M_AXI_ARVALID;
  assign io_M_AXI_1_WDATA = MAGToAXI4Bridge_1_io_M_AXI_WDATA;
  assign io_M_AXI_1_WSTRB = MAGToAXI4Bridge_1_io_M_AXI_WSTRB;
  assign io_M_AXI_1_WVALID = MAGToAXI4Bridge_1_io_M_AXI_WVALID;
  assign io_M_AXI_1_RREADY = MAGToAXI4Bridge_1_io_M_AXI_RREADY;
  assign io_M_AXI_1_BREADY = MAGToAXI4Bridge_1_io_M_AXI_BREADY;
  assign io_M_AXI_2_AWID = MAGToAXI4Bridge_2_io_M_AXI_AWID;
  assign io_M_AXI_2_AWADDR = MAGToAXI4Bridge_2_io_M_AXI_AWADDR;
  assign io_M_AXI_2_AWLEN = MAGToAXI4Bridge_2_io_M_AXI_AWLEN;
  assign io_M_AXI_2_AWVALID = MAGToAXI4Bridge_2_io_M_AXI_AWVALID;
  assign io_M_AXI_2_ARID = MAGToAXI4Bridge_2_io_M_AXI_ARID;
  assign io_M_AXI_2_ARADDR = MAGToAXI4Bridge_2_io_M_AXI_ARADDR;
  assign io_M_AXI_2_ARLEN = MAGToAXI4Bridge_2_io_M_AXI_ARLEN;
  assign io_M_AXI_2_ARVALID = MAGToAXI4Bridge_2_io_M_AXI_ARVALID;
  assign io_M_AXI_2_WDATA = MAGToAXI4Bridge_2_io_M_AXI_WDATA;
  assign io_M_AXI_2_WSTRB = MAGToAXI4Bridge_2_io_M_AXI_WSTRB;
  assign io_M_AXI_2_WVALID = MAGToAXI4Bridge_2_io_M_AXI_WVALID;
  assign io_M_AXI_2_RREADY = MAGToAXI4Bridge_2_io_M_AXI_RREADY;
  assign io_M_AXI_2_BREADY = MAGToAXI4Bridge_2_io_M_AXI_BREADY;
  assign io_M_AXI_3_AWID = MAGToAXI4Bridge_3_io_M_AXI_AWID;
  assign io_M_AXI_3_AWADDR = MAGToAXI4Bridge_3_io_M_AXI_AWADDR;
  assign io_M_AXI_3_AWLEN = MAGToAXI4Bridge_3_io_M_AXI_AWLEN;
  assign io_M_AXI_3_AWVALID = MAGToAXI4Bridge_3_io_M_AXI_AWVALID;
  assign io_M_AXI_3_ARID = MAGToAXI4Bridge_3_io_M_AXI_ARID;
  assign io_M_AXI_3_ARADDR = MAGToAXI4Bridge_3_io_M_AXI_ARADDR;
  assign io_M_AXI_3_ARLEN = MAGToAXI4Bridge_3_io_M_AXI_ARLEN;
  assign io_M_AXI_3_ARVALID = MAGToAXI4Bridge_3_io_M_AXI_ARVALID;
  assign io_M_AXI_3_WDATA = MAGToAXI4Bridge_3_io_M_AXI_WDATA;
  assign io_M_AXI_3_WSTRB = MAGToAXI4Bridge_3_io_M_AXI_WSTRB;
  assign io_M_AXI_3_WVALID = MAGToAXI4Bridge_3_io_M_AXI_WVALID;
  assign io_M_AXI_3_RREADY = MAGToAXI4Bridge_3_io_M_AXI_RREADY;
  assign io_M_AXI_3_BREADY = MAGToAXI4Bridge_3_io_M_AXI_BREADY;
  assign io_enable = fringeCommon_io_enable;
  assign io_reset = fringeCommon_io_reset;
  assign io_argIns_0 = fringeCommon_io_argIns_0;
  assign io_argIns_1 = fringeCommon_io_argIns_1;
  assign io_argIns_2 = fringeCommon_io_argIns_2;
  assign io_memStreams_loads_3_cmd_ready = fringeCommon_io_memStreams_loads_3_cmd_ready;
  assign io_memStreams_loads_3_rdata_valid = fringeCommon_io_memStreams_loads_3_rdata_valid;
  assign io_memStreams_loads_3_rdata_bits_0 = fringeCommon_io_memStreams_loads_3_rdata_bits_0;
  assign io_memStreams_loads_2_cmd_ready = fringeCommon_io_memStreams_loads_2_cmd_ready;
  assign io_memStreams_loads_2_rdata_valid = fringeCommon_io_memStreams_loads_2_rdata_valid;
  assign io_memStreams_loads_2_rdata_bits_0 = fringeCommon_io_memStreams_loads_2_rdata_bits_0;
  assign io_memStreams_loads_1_cmd_ready = fringeCommon_io_memStreams_loads_1_cmd_ready;
  assign io_memStreams_loads_1_rdata_valid = fringeCommon_io_memStreams_loads_1_rdata_valid;
  assign io_memStreams_loads_1_rdata_bits_0 = fringeCommon_io_memStreams_loads_1_rdata_bits_0;
  assign io_memStreams_loads_0_cmd_ready = fringeCommon_io_memStreams_loads_0_cmd_ready;
  assign io_memStreams_loads_0_rdata_valid = fringeCommon_io_memStreams_loads_0_rdata_valid;
  assign io_memStreams_loads_0_rdata_bits_0 = fringeCommon_io_memStreams_loads_0_rdata_bits_0;
  assign fringeCommon_io_raddr = AXI4LiteToRFBridge_io_raddr;
  assign fringeCommon_io_wen = AXI4LiteToRFBridge_io_wen;
  assign fringeCommon_io_waddr = AXI4LiteToRFBridge_io_waddr;
  assign fringeCommon_io_wdata = {{32'd0}, AXI4LiteToRFBridge_io_wdata};
  assign fringeCommon_io_done = io_done;
  assign fringeCommon_io_argOuts_0_valid = io_argOuts_0_valid;
  assign fringeCommon_io_argOuts_0_bits = io_argOuts_0_bits;
  assign fringeCommon_io_memStreams_loads_3_cmd_valid = io_memStreams_loads_3_cmd_valid;
  assign fringeCommon_io_memStreams_loads_3_cmd_bits_addr = io_memStreams_loads_3_cmd_bits_addr;
  assign fringeCommon_io_memStreams_loads_3_cmd_bits_isWr = io_memStreams_loads_3_cmd_bits_isWr;
  assign fringeCommon_io_memStreams_loads_3_cmd_bits_size = io_memStreams_loads_3_cmd_bits_size;
  assign fringeCommon_io_memStreams_loads_3_rdata_ready = io_memStreams_loads_3_rdata_ready;
  assign fringeCommon_io_memStreams_loads_2_cmd_valid = io_memStreams_loads_2_cmd_valid;
  assign fringeCommon_io_memStreams_loads_2_cmd_bits_addr = io_memStreams_loads_2_cmd_bits_addr;
  assign fringeCommon_io_memStreams_loads_2_cmd_bits_isWr = io_memStreams_loads_2_cmd_bits_isWr;
  assign fringeCommon_io_memStreams_loads_2_cmd_bits_size = io_memStreams_loads_2_cmd_bits_size;
  assign fringeCommon_io_memStreams_loads_2_rdata_ready = io_memStreams_loads_2_rdata_ready;
  assign fringeCommon_io_memStreams_loads_1_cmd_valid = io_memStreams_loads_1_cmd_valid;
  assign fringeCommon_io_memStreams_loads_1_cmd_bits_addr = io_memStreams_loads_1_cmd_bits_addr;
  assign fringeCommon_io_memStreams_loads_1_cmd_bits_isWr = io_memStreams_loads_1_cmd_bits_isWr;
  assign fringeCommon_io_memStreams_loads_1_cmd_bits_size = io_memStreams_loads_1_cmd_bits_size;
  assign fringeCommon_io_memStreams_loads_1_rdata_ready = io_memStreams_loads_1_rdata_ready;
  assign fringeCommon_io_memStreams_loads_0_cmd_valid = io_memStreams_loads_0_cmd_valid;
  assign fringeCommon_io_memStreams_loads_0_cmd_bits_addr = io_memStreams_loads_0_cmd_bits_addr;
  assign fringeCommon_io_memStreams_loads_0_cmd_bits_isWr = io_memStreams_loads_0_cmd_bits_isWr;
  assign fringeCommon_io_memStreams_loads_0_cmd_bits_size = io_memStreams_loads_0_cmd_bits_size;
  assign fringeCommon_io_memStreams_loads_0_rdata_ready = io_memStreams_loads_0_rdata_ready;
  assign fringeCommon_io_dram_0_cmd_ready = MAGToAXI4Bridge_io_in_cmd_ready;
  assign fringeCommon_io_dram_0_wdata_ready = MAGToAXI4Bridge_io_in_wdata_ready;
  assign fringeCommon_io_dram_0_rresp_valid = MAGToAXI4Bridge_io_in_rresp_valid;
  assign fringeCommon_io_dram_0_rresp_bits_rdata_0 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_0;
  assign fringeCommon_io_dram_0_rresp_bits_rdata_1 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_1;
  assign fringeCommon_io_dram_0_rresp_bits_rdata_2 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_2;
  assign fringeCommon_io_dram_0_rresp_bits_rdata_3 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_3;
  assign fringeCommon_io_dram_0_rresp_bits_rdata_4 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_4;
  assign fringeCommon_io_dram_0_rresp_bits_rdata_5 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_5;
  assign fringeCommon_io_dram_0_rresp_bits_rdata_6 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_6;
  assign fringeCommon_io_dram_0_rresp_bits_rdata_7 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_7;
  assign fringeCommon_io_dram_0_rresp_bits_rdata_8 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_8;
  assign fringeCommon_io_dram_0_rresp_bits_rdata_9 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_9;
  assign fringeCommon_io_dram_0_rresp_bits_rdata_10 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_10;
  assign fringeCommon_io_dram_0_rresp_bits_rdata_11 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_11;
  assign fringeCommon_io_dram_0_rresp_bits_rdata_12 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_12;
  assign fringeCommon_io_dram_0_rresp_bits_rdata_13 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_13;
  assign fringeCommon_io_dram_0_rresp_bits_rdata_14 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_14;
  assign fringeCommon_io_dram_0_rresp_bits_rdata_15 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_15;
  assign fringeCommon_io_dram_0_rresp_bits_tag_streamId = MAGToAXI4Bridge_io_in_rresp_bits_tag_streamId;
  assign fringeCommon_io_dram_0_wresp_valid = MAGToAXI4Bridge_io_in_wresp_valid;
  assign fringeCommon_io_dram_0_wresp_bits_tag_streamId = MAGToAXI4Bridge_io_in_wresp_bits_tag_streamId;
  assign fringeCommon_io_dram_1_cmd_ready = MAGToAXI4Bridge_1_io_in_cmd_ready;
  assign fringeCommon_io_dram_1_wdata_ready = MAGToAXI4Bridge_1_io_in_wdata_ready;
  assign fringeCommon_io_dram_1_rresp_valid = MAGToAXI4Bridge_1_io_in_rresp_valid;
  assign fringeCommon_io_dram_1_rresp_bits_rdata_0 = MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_0;
  assign fringeCommon_io_dram_1_rresp_bits_rdata_1 = MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_1;
  assign fringeCommon_io_dram_1_rresp_bits_rdata_2 = MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_2;
  assign fringeCommon_io_dram_1_rresp_bits_rdata_3 = MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_3;
  assign fringeCommon_io_dram_1_rresp_bits_rdata_4 = MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_4;
  assign fringeCommon_io_dram_1_rresp_bits_rdata_5 = MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_5;
  assign fringeCommon_io_dram_1_rresp_bits_rdata_6 = MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_6;
  assign fringeCommon_io_dram_1_rresp_bits_rdata_7 = MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_7;
  assign fringeCommon_io_dram_1_rresp_bits_rdata_8 = MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_8;
  assign fringeCommon_io_dram_1_rresp_bits_rdata_9 = MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_9;
  assign fringeCommon_io_dram_1_rresp_bits_rdata_10 = MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_10;
  assign fringeCommon_io_dram_1_rresp_bits_rdata_11 = MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_11;
  assign fringeCommon_io_dram_1_rresp_bits_rdata_12 = MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_12;
  assign fringeCommon_io_dram_1_rresp_bits_rdata_13 = MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_13;
  assign fringeCommon_io_dram_1_rresp_bits_rdata_14 = MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_14;
  assign fringeCommon_io_dram_1_rresp_bits_rdata_15 = MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_15;
  assign fringeCommon_io_dram_1_rresp_bits_tag_streamId = MAGToAXI4Bridge_1_io_in_rresp_bits_tag_streamId;
  assign fringeCommon_io_dram_1_wresp_valid = MAGToAXI4Bridge_1_io_in_wresp_valid;
  assign fringeCommon_io_dram_1_wresp_bits_tag_streamId = MAGToAXI4Bridge_1_io_in_wresp_bits_tag_streamId;
  assign fringeCommon_io_dram_2_cmd_ready = MAGToAXI4Bridge_2_io_in_cmd_ready;
  assign fringeCommon_io_dram_2_wdata_ready = MAGToAXI4Bridge_2_io_in_wdata_ready;
  assign fringeCommon_io_dram_2_rresp_valid = MAGToAXI4Bridge_2_io_in_rresp_valid;
  assign fringeCommon_io_dram_2_rresp_bits_rdata_0 = MAGToAXI4Bridge_2_io_in_rresp_bits_rdata_0;
  assign fringeCommon_io_dram_2_rresp_bits_rdata_1 = MAGToAXI4Bridge_2_io_in_rresp_bits_rdata_1;
  assign fringeCommon_io_dram_2_rresp_bits_rdata_2 = MAGToAXI4Bridge_2_io_in_rresp_bits_rdata_2;
  assign fringeCommon_io_dram_2_rresp_bits_rdata_3 = MAGToAXI4Bridge_2_io_in_rresp_bits_rdata_3;
  assign fringeCommon_io_dram_2_rresp_bits_rdata_4 = MAGToAXI4Bridge_2_io_in_rresp_bits_rdata_4;
  assign fringeCommon_io_dram_2_rresp_bits_rdata_5 = MAGToAXI4Bridge_2_io_in_rresp_bits_rdata_5;
  assign fringeCommon_io_dram_2_rresp_bits_rdata_6 = MAGToAXI4Bridge_2_io_in_rresp_bits_rdata_6;
  assign fringeCommon_io_dram_2_rresp_bits_rdata_7 = MAGToAXI4Bridge_2_io_in_rresp_bits_rdata_7;
  assign fringeCommon_io_dram_2_rresp_bits_rdata_8 = MAGToAXI4Bridge_2_io_in_rresp_bits_rdata_8;
  assign fringeCommon_io_dram_2_rresp_bits_rdata_9 = MAGToAXI4Bridge_2_io_in_rresp_bits_rdata_9;
  assign fringeCommon_io_dram_2_rresp_bits_rdata_10 = MAGToAXI4Bridge_2_io_in_rresp_bits_rdata_10;
  assign fringeCommon_io_dram_2_rresp_bits_rdata_11 = MAGToAXI4Bridge_2_io_in_rresp_bits_rdata_11;
  assign fringeCommon_io_dram_2_rresp_bits_rdata_12 = MAGToAXI4Bridge_2_io_in_rresp_bits_rdata_12;
  assign fringeCommon_io_dram_2_rresp_bits_rdata_13 = MAGToAXI4Bridge_2_io_in_rresp_bits_rdata_13;
  assign fringeCommon_io_dram_2_rresp_bits_rdata_14 = MAGToAXI4Bridge_2_io_in_rresp_bits_rdata_14;
  assign fringeCommon_io_dram_2_rresp_bits_rdata_15 = MAGToAXI4Bridge_2_io_in_rresp_bits_rdata_15;
  assign fringeCommon_io_dram_2_rresp_bits_tag_streamId = MAGToAXI4Bridge_2_io_in_rresp_bits_tag_streamId;
  assign fringeCommon_io_dram_2_wresp_valid = MAGToAXI4Bridge_2_io_in_wresp_valid;
  assign fringeCommon_io_dram_2_wresp_bits_tag_streamId = MAGToAXI4Bridge_2_io_in_wresp_bits_tag_streamId;
  assign fringeCommon_io_dram_3_cmd_ready = MAGToAXI4Bridge_3_io_in_cmd_ready;
  assign fringeCommon_io_dram_3_wdata_ready = MAGToAXI4Bridge_3_io_in_wdata_ready;
  assign fringeCommon_io_dram_3_rresp_valid = MAGToAXI4Bridge_3_io_in_rresp_valid;
  assign fringeCommon_io_dram_3_rresp_bits_rdata_0 = MAGToAXI4Bridge_3_io_in_rresp_bits_rdata_0;
  assign fringeCommon_io_dram_3_rresp_bits_rdata_1 = MAGToAXI4Bridge_3_io_in_rresp_bits_rdata_1;
  assign fringeCommon_io_dram_3_rresp_bits_rdata_2 = MAGToAXI4Bridge_3_io_in_rresp_bits_rdata_2;
  assign fringeCommon_io_dram_3_rresp_bits_rdata_3 = MAGToAXI4Bridge_3_io_in_rresp_bits_rdata_3;
  assign fringeCommon_io_dram_3_rresp_bits_rdata_4 = MAGToAXI4Bridge_3_io_in_rresp_bits_rdata_4;
  assign fringeCommon_io_dram_3_rresp_bits_rdata_5 = MAGToAXI4Bridge_3_io_in_rresp_bits_rdata_5;
  assign fringeCommon_io_dram_3_rresp_bits_rdata_6 = MAGToAXI4Bridge_3_io_in_rresp_bits_rdata_6;
  assign fringeCommon_io_dram_3_rresp_bits_rdata_7 = MAGToAXI4Bridge_3_io_in_rresp_bits_rdata_7;
  assign fringeCommon_io_dram_3_rresp_bits_rdata_8 = MAGToAXI4Bridge_3_io_in_rresp_bits_rdata_8;
  assign fringeCommon_io_dram_3_rresp_bits_rdata_9 = MAGToAXI4Bridge_3_io_in_rresp_bits_rdata_9;
  assign fringeCommon_io_dram_3_rresp_bits_rdata_10 = MAGToAXI4Bridge_3_io_in_rresp_bits_rdata_10;
  assign fringeCommon_io_dram_3_rresp_bits_rdata_11 = MAGToAXI4Bridge_3_io_in_rresp_bits_rdata_11;
  assign fringeCommon_io_dram_3_rresp_bits_rdata_12 = MAGToAXI4Bridge_3_io_in_rresp_bits_rdata_12;
  assign fringeCommon_io_dram_3_rresp_bits_rdata_13 = MAGToAXI4Bridge_3_io_in_rresp_bits_rdata_13;
  assign fringeCommon_io_dram_3_rresp_bits_rdata_14 = MAGToAXI4Bridge_3_io_in_rresp_bits_rdata_14;
  assign fringeCommon_io_dram_3_rresp_bits_rdata_15 = MAGToAXI4Bridge_3_io_in_rresp_bits_rdata_15;
  assign fringeCommon_io_dram_3_rresp_bits_tag_streamId = MAGToAXI4Bridge_3_io_in_rresp_bits_tag_streamId;
  assign fringeCommon_io_dram_3_wresp_valid = MAGToAXI4Bridge_3_io_in_wresp_valid;
  assign fringeCommon_io_dram_3_wresp_bits_tag_streamId = MAGToAXI4Bridge_3_io_in_wresp_bits_tag_streamId;
  assign fringeCommon_io_TOP_AXI_AWADDR = {{32'd0}, io_TOP_AXI_AWADDR};
  assign fringeCommon_io_TOP_AXI_AWLEN = io_TOP_AXI_AWLEN;
  assign fringeCommon_io_TOP_AXI_AWVALID = io_TOP_AXI_AWVALID;
  assign fringeCommon_io_TOP_AXI_AWREADY = io_TOP_AXI_AWREADY;
  assign fringeCommon_io_TOP_AXI_ARID = io_TOP_AXI_ARID;
  assign fringeCommon_io_TOP_AXI_ARADDR = {{32'd0}, io_TOP_AXI_ARADDR};
  assign fringeCommon_io_TOP_AXI_ARLEN = io_TOP_AXI_ARLEN;
  assign fringeCommon_io_TOP_AXI_ARSIZE = io_TOP_AXI_ARSIZE;
  assign fringeCommon_io_TOP_AXI_ARBURST = io_TOP_AXI_ARBURST;
  assign fringeCommon_io_TOP_AXI_ARVALID = io_TOP_AXI_ARVALID;
  assign fringeCommon_io_TOP_AXI_ARREADY = io_TOP_AXI_ARREADY;
  assign fringeCommon_io_TOP_AXI_WDATA = {{480'd0}, io_TOP_AXI_WDATA};
  assign fringeCommon_io_TOP_AXI_WSTRB = io_TOP_AXI_WSTRB;
  assign fringeCommon_io_TOP_AXI_WVALID = io_TOP_AXI_WVALID;
  assign fringeCommon_io_TOP_AXI_WREADY = io_TOP_AXI_WREADY;
  assign fringeCommon_io_TOP_AXI_RVALID = io_TOP_AXI_RVALID;
  assign fringeCommon_io_TOP_AXI_RREADY = io_TOP_AXI_RREADY;
  assign fringeCommon_io_TOP_AXI_BVALID = io_TOP_AXI_BVALID;
  assign fringeCommon_io_TOP_AXI_BREADY = io_TOP_AXI_BREADY;
  assign fringeCommon_io_DWIDTH_AXI_AWADDR = {{32'd0}, io_DWIDTH_AXI_AWADDR};
  assign fringeCommon_io_DWIDTH_AXI_AWLEN = io_DWIDTH_AXI_AWLEN;
  assign fringeCommon_io_DWIDTH_AXI_AWVALID = io_DWIDTH_AXI_AWVALID;
  assign fringeCommon_io_DWIDTH_AXI_AWREADY = io_DWIDTH_AXI_AWREADY;
  assign fringeCommon_io_DWIDTH_AXI_ARADDR = {{32'd0}, io_DWIDTH_AXI_ARADDR};
  assign fringeCommon_io_DWIDTH_AXI_ARLEN = io_DWIDTH_AXI_ARLEN;
  assign fringeCommon_io_DWIDTH_AXI_ARSIZE = io_DWIDTH_AXI_ARSIZE;
  assign fringeCommon_io_DWIDTH_AXI_ARBURST = io_DWIDTH_AXI_ARBURST;
  assign fringeCommon_io_DWIDTH_AXI_ARVALID = io_DWIDTH_AXI_ARVALID;
  assign fringeCommon_io_DWIDTH_AXI_ARREADY = io_DWIDTH_AXI_ARREADY;
  assign fringeCommon_io_DWIDTH_AXI_WDATA = {{480'd0}, io_DWIDTH_AXI_WDATA};
  assign fringeCommon_io_DWIDTH_AXI_WSTRB = io_DWIDTH_AXI_WSTRB;
  assign fringeCommon_io_DWIDTH_AXI_WVALID = io_DWIDTH_AXI_WVALID;
  assign fringeCommon_io_DWIDTH_AXI_WREADY = io_DWIDTH_AXI_WREADY;
  assign fringeCommon_io_DWIDTH_AXI_RVALID = io_DWIDTH_AXI_RVALID;
  assign fringeCommon_io_DWIDTH_AXI_RREADY = io_DWIDTH_AXI_RREADY;
  assign fringeCommon_io_DWIDTH_AXI_BVALID = io_DWIDTH_AXI_BVALID;
  assign fringeCommon_io_DWIDTH_AXI_BREADY = io_DWIDTH_AXI_BREADY;
  assign fringeCommon_clock = clock;
  assign fringeCommon_reset = reset;
  assign AXI4LiteToRFBridge_io_S_AXI_AWADDR = io_S_AXI_AWADDR;
  assign AXI4LiteToRFBridge_io_S_AXI_AWPROT = io_S_AXI_AWPROT;
  assign AXI4LiteToRFBridge_io_S_AXI_AWVALID = io_S_AXI_AWVALID;
  assign AXI4LiteToRFBridge_io_S_AXI_ARADDR = io_S_AXI_ARADDR;
  assign AXI4LiteToRFBridge_io_S_AXI_ARPROT = io_S_AXI_ARPROT;
  assign AXI4LiteToRFBridge_io_S_AXI_ARVALID = io_S_AXI_ARVALID;
  assign AXI4LiteToRFBridge_io_S_AXI_WDATA = io_S_AXI_WDATA;
  assign AXI4LiteToRFBridge_io_S_AXI_WSTRB = io_S_AXI_WSTRB;
  assign AXI4LiteToRFBridge_io_S_AXI_WVALID = io_S_AXI_WVALID;
  assign AXI4LiteToRFBridge_io_S_AXI_RREADY = io_S_AXI_RREADY;
  assign AXI4LiteToRFBridge_io_S_AXI_BREADY = io_S_AXI_BREADY;
  assign AXI4LiteToRFBridge_io_rdata = fringeCommon_io_rdata[31:0];
  assign AXI4LiteToRFBridge_clock = clock;
  assign AXI4LiteToRFBridge_reset = reset;
  assign MAGToAXI4Bridge_io_in_cmd_valid = fringeCommon_io_dram_0_cmd_valid;
  assign MAGToAXI4Bridge_io_in_cmd_bits_addr = fringeCommon_io_dram_0_cmd_bits_addr;
  assign MAGToAXI4Bridge_io_in_cmd_bits_size = fringeCommon_io_dram_0_cmd_bits_size;
  assign MAGToAXI4Bridge_io_in_cmd_bits_isWr = fringeCommon_io_dram_0_cmd_bits_isWr;
  assign MAGToAXI4Bridge_io_in_cmd_bits_tag_uid = fringeCommon_io_dram_0_cmd_bits_tag_uid;
  assign MAGToAXI4Bridge_io_in_cmd_bits_tag_streamId = fringeCommon_io_dram_0_cmd_bits_tag_streamId;
  assign MAGToAXI4Bridge_io_in_wdata_valid = fringeCommon_io_dram_0_wdata_valid;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_0_wdata_bits_wdata_0;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_0_wdata_bits_wdata_1;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_0_wdata_bits_wdata_2;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_0_wdata_bits_wdata_3;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_0_wdata_bits_wdata_4;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_0_wdata_bits_wdata_5;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_0_wdata_bits_wdata_6;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_0_wdata_bits_wdata_7;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_0_wdata_bits_wdata_8;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_0_wdata_bits_wdata_9;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_0_wdata_bits_wdata_10;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_0_wdata_bits_wdata_11;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_0_wdata_bits_wdata_12;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_0_wdata_bits_wdata_13;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_0_wdata_bits_wdata_14;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_0_wdata_bits_wdata_15;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_0_wdata_bits_wstrb_0;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_0_wdata_bits_wstrb_1;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_0_wdata_bits_wstrb_2;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_0_wdata_bits_wstrb_3;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_0_wdata_bits_wstrb_4;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_0_wdata_bits_wstrb_5;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_0_wdata_bits_wstrb_6;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_0_wdata_bits_wstrb_7;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_0_wdata_bits_wstrb_8;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_0_wdata_bits_wstrb_9;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_0_wdata_bits_wstrb_10;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_0_wdata_bits_wstrb_11;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_0_wdata_bits_wstrb_12;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_0_wdata_bits_wstrb_13;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_0_wdata_bits_wstrb_14;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_0_wdata_bits_wstrb_15;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_0_wdata_bits_wstrb_16;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_0_wdata_bits_wstrb_17;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_0_wdata_bits_wstrb_18;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_0_wdata_bits_wstrb_19;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_0_wdata_bits_wstrb_20;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_0_wdata_bits_wstrb_21;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_0_wdata_bits_wstrb_22;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_0_wdata_bits_wstrb_23;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_0_wdata_bits_wstrb_24;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_0_wdata_bits_wstrb_25;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_0_wdata_bits_wstrb_26;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_0_wdata_bits_wstrb_27;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_0_wdata_bits_wstrb_28;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_0_wdata_bits_wstrb_29;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_0_wdata_bits_wstrb_30;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_0_wdata_bits_wstrb_31;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_0_wdata_bits_wstrb_32;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_0_wdata_bits_wstrb_33;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_0_wdata_bits_wstrb_34;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_0_wdata_bits_wstrb_35;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_0_wdata_bits_wstrb_36;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_0_wdata_bits_wstrb_37;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_0_wdata_bits_wstrb_38;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_0_wdata_bits_wstrb_39;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_0_wdata_bits_wstrb_40;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_0_wdata_bits_wstrb_41;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_0_wdata_bits_wstrb_42;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_0_wdata_bits_wstrb_43;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_0_wdata_bits_wstrb_44;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_0_wdata_bits_wstrb_45;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_0_wdata_bits_wstrb_46;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_0_wdata_bits_wstrb_47;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_0_wdata_bits_wstrb_48;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_0_wdata_bits_wstrb_49;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_0_wdata_bits_wstrb_50;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_0_wdata_bits_wstrb_51;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_0_wdata_bits_wstrb_52;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_0_wdata_bits_wstrb_53;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_0_wdata_bits_wstrb_54;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_0_wdata_bits_wstrb_55;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_0_wdata_bits_wstrb_56;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_0_wdata_bits_wstrb_57;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_0_wdata_bits_wstrb_58;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_0_wdata_bits_wstrb_59;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_0_wdata_bits_wstrb_60;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_0_wdata_bits_wstrb_61;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_0_wdata_bits_wstrb_62;
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_0_wdata_bits_wstrb_63;
  assign MAGToAXI4Bridge_io_in_rresp_ready = fringeCommon_io_dram_0_rresp_ready;
  assign MAGToAXI4Bridge_io_in_wresp_ready = fringeCommon_io_dram_0_wresp_ready;
  assign MAGToAXI4Bridge_io_M_AXI_AWREADY = io_M_AXI_0_AWREADY;
  assign MAGToAXI4Bridge_io_M_AXI_ARREADY = io_M_AXI_0_ARREADY;
  assign MAGToAXI4Bridge_io_M_AXI_WREADY = io_M_AXI_0_WREADY;
  assign MAGToAXI4Bridge_io_M_AXI_RID = io_M_AXI_0_RID;
  assign MAGToAXI4Bridge_io_M_AXI_RDATA = io_M_AXI_0_RDATA;
  assign MAGToAXI4Bridge_io_M_AXI_RVALID = io_M_AXI_0_RVALID;
  assign MAGToAXI4Bridge_io_M_AXI_BID = io_M_AXI_0_BID;
  assign MAGToAXI4Bridge_io_M_AXI_BVALID = io_M_AXI_0_BVALID;
  assign MAGToAXI4Bridge_1_io_in_cmd_valid = fringeCommon_io_dram_1_cmd_valid;
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_addr = fringeCommon_io_dram_1_cmd_bits_addr;
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_size = fringeCommon_io_dram_1_cmd_bits_size;
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_isWr = fringeCommon_io_dram_1_cmd_bits_isWr;
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_tag_uid = fringeCommon_io_dram_1_cmd_bits_tag_uid;
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_tag_streamId = fringeCommon_io_dram_1_cmd_bits_tag_streamId;
  assign MAGToAXI4Bridge_1_io_in_wdata_valid = fringeCommon_io_dram_1_wdata_valid;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_1_wdata_bits_wdata_0;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_1_wdata_bits_wdata_1;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_1_wdata_bits_wdata_2;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_1_wdata_bits_wdata_3;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_1_wdata_bits_wdata_4;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_1_wdata_bits_wdata_5;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_1_wdata_bits_wdata_6;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_1_wdata_bits_wdata_7;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_1_wdata_bits_wdata_8;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_1_wdata_bits_wdata_9;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_1_wdata_bits_wdata_10;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_1_wdata_bits_wdata_11;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_1_wdata_bits_wdata_12;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_1_wdata_bits_wdata_13;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_1_wdata_bits_wdata_14;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_1_wdata_bits_wdata_15;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_1_wdata_bits_wstrb_0;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_1_wdata_bits_wstrb_1;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_1_wdata_bits_wstrb_2;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_1_wdata_bits_wstrb_3;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_1_wdata_bits_wstrb_4;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_1_wdata_bits_wstrb_5;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_1_wdata_bits_wstrb_6;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_1_wdata_bits_wstrb_7;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_1_wdata_bits_wstrb_8;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_1_wdata_bits_wstrb_9;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_1_wdata_bits_wstrb_10;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_1_wdata_bits_wstrb_11;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_1_wdata_bits_wstrb_12;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_1_wdata_bits_wstrb_13;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_1_wdata_bits_wstrb_14;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_1_wdata_bits_wstrb_15;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_1_wdata_bits_wstrb_16;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_1_wdata_bits_wstrb_17;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_1_wdata_bits_wstrb_18;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_1_wdata_bits_wstrb_19;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_1_wdata_bits_wstrb_20;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_1_wdata_bits_wstrb_21;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_1_wdata_bits_wstrb_22;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_1_wdata_bits_wstrb_23;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_1_wdata_bits_wstrb_24;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_1_wdata_bits_wstrb_25;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_1_wdata_bits_wstrb_26;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_1_wdata_bits_wstrb_27;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_1_wdata_bits_wstrb_28;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_1_wdata_bits_wstrb_29;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_1_wdata_bits_wstrb_30;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_1_wdata_bits_wstrb_31;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_1_wdata_bits_wstrb_32;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_1_wdata_bits_wstrb_33;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_1_wdata_bits_wstrb_34;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_1_wdata_bits_wstrb_35;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_1_wdata_bits_wstrb_36;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_1_wdata_bits_wstrb_37;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_1_wdata_bits_wstrb_38;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_1_wdata_bits_wstrb_39;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_1_wdata_bits_wstrb_40;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_1_wdata_bits_wstrb_41;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_1_wdata_bits_wstrb_42;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_1_wdata_bits_wstrb_43;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_1_wdata_bits_wstrb_44;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_1_wdata_bits_wstrb_45;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_1_wdata_bits_wstrb_46;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_1_wdata_bits_wstrb_47;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_1_wdata_bits_wstrb_48;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_1_wdata_bits_wstrb_49;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_1_wdata_bits_wstrb_50;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_1_wdata_bits_wstrb_51;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_1_wdata_bits_wstrb_52;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_1_wdata_bits_wstrb_53;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_1_wdata_bits_wstrb_54;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_1_wdata_bits_wstrb_55;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_1_wdata_bits_wstrb_56;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_1_wdata_bits_wstrb_57;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_1_wdata_bits_wstrb_58;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_1_wdata_bits_wstrb_59;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_1_wdata_bits_wstrb_60;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_1_wdata_bits_wstrb_61;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_1_wdata_bits_wstrb_62;
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_1_wdata_bits_wstrb_63;
  assign MAGToAXI4Bridge_1_io_in_rresp_ready = fringeCommon_io_dram_1_rresp_ready;
  assign MAGToAXI4Bridge_1_io_in_wresp_ready = fringeCommon_io_dram_1_wresp_ready;
  assign MAGToAXI4Bridge_1_io_M_AXI_AWREADY = io_M_AXI_1_AWREADY;
  assign MAGToAXI4Bridge_1_io_M_AXI_ARREADY = io_M_AXI_1_ARREADY;
  assign MAGToAXI4Bridge_1_io_M_AXI_WREADY = io_M_AXI_1_WREADY;
  assign MAGToAXI4Bridge_1_io_M_AXI_RID = io_M_AXI_1_RID;
  assign MAGToAXI4Bridge_1_io_M_AXI_RDATA = io_M_AXI_1_RDATA;
  assign MAGToAXI4Bridge_1_io_M_AXI_RVALID = io_M_AXI_1_RVALID;
  assign MAGToAXI4Bridge_1_io_M_AXI_BID = io_M_AXI_1_BID;
  assign MAGToAXI4Bridge_1_io_M_AXI_BVALID = io_M_AXI_1_BVALID;
  assign MAGToAXI4Bridge_2_io_in_cmd_valid = fringeCommon_io_dram_2_cmd_valid;
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_addr = fringeCommon_io_dram_2_cmd_bits_addr;
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_size = fringeCommon_io_dram_2_cmd_bits_size;
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_isWr = fringeCommon_io_dram_2_cmd_bits_isWr;
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_tag_uid = fringeCommon_io_dram_2_cmd_bits_tag_uid;
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_tag_streamId = fringeCommon_io_dram_2_cmd_bits_tag_streamId;
  assign MAGToAXI4Bridge_2_io_in_wdata_valid = fringeCommon_io_dram_2_wdata_valid;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_2_wdata_bits_wdata_0;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_2_wdata_bits_wdata_1;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_2_wdata_bits_wdata_2;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_2_wdata_bits_wdata_3;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_2_wdata_bits_wdata_4;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_2_wdata_bits_wdata_5;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_2_wdata_bits_wdata_6;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_2_wdata_bits_wdata_7;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_2_wdata_bits_wdata_8;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_2_wdata_bits_wdata_9;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_2_wdata_bits_wdata_10;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_2_wdata_bits_wdata_11;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_2_wdata_bits_wdata_12;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_2_wdata_bits_wdata_13;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_2_wdata_bits_wdata_14;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_2_wdata_bits_wdata_15;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_2_wdata_bits_wstrb_0;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_2_wdata_bits_wstrb_1;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_2_wdata_bits_wstrb_2;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_2_wdata_bits_wstrb_3;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_2_wdata_bits_wstrb_4;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_2_wdata_bits_wstrb_5;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_2_wdata_bits_wstrb_6;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_2_wdata_bits_wstrb_7;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_2_wdata_bits_wstrb_8;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_2_wdata_bits_wstrb_9;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_2_wdata_bits_wstrb_10;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_2_wdata_bits_wstrb_11;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_2_wdata_bits_wstrb_12;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_2_wdata_bits_wstrb_13;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_2_wdata_bits_wstrb_14;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_2_wdata_bits_wstrb_15;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_2_wdata_bits_wstrb_16;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_2_wdata_bits_wstrb_17;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_2_wdata_bits_wstrb_18;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_2_wdata_bits_wstrb_19;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_2_wdata_bits_wstrb_20;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_2_wdata_bits_wstrb_21;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_2_wdata_bits_wstrb_22;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_2_wdata_bits_wstrb_23;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_2_wdata_bits_wstrb_24;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_2_wdata_bits_wstrb_25;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_2_wdata_bits_wstrb_26;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_2_wdata_bits_wstrb_27;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_2_wdata_bits_wstrb_28;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_2_wdata_bits_wstrb_29;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_2_wdata_bits_wstrb_30;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_2_wdata_bits_wstrb_31;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_2_wdata_bits_wstrb_32;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_2_wdata_bits_wstrb_33;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_2_wdata_bits_wstrb_34;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_2_wdata_bits_wstrb_35;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_2_wdata_bits_wstrb_36;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_2_wdata_bits_wstrb_37;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_2_wdata_bits_wstrb_38;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_2_wdata_bits_wstrb_39;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_2_wdata_bits_wstrb_40;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_2_wdata_bits_wstrb_41;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_2_wdata_bits_wstrb_42;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_2_wdata_bits_wstrb_43;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_2_wdata_bits_wstrb_44;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_2_wdata_bits_wstrb_45;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_2_wdata_bits_wstrb_46;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_2_wdata_bits_wstrb_47;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_2_wdata_bits_wstrb_48;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_2_wdata_bits_wstrb_49;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_2_wdata_bits_wstrb_50;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_2_wdata_bits_wstrb_51;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_2_wdata_bits_wstrb_52;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_2_wdata_bits_wstrb_53;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_2_wdata_bits_wstrb_54;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_2_wdata_bits_wstrb_55;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_2_wdata_bits_wstrb_56;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_2_wdata_bits_wstrb_57;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_2_wdata_bits_wstrb_58;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_2_wdata_bits_wstrb_59;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_2_wdata_bits_wstrb_60;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_2_wdata_bits_wstrb_61;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_2_wdata_bits_wstrb_62;
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_2_wdata_bits_wstrb_63;
  assign MAGToAXI4Bridge_2_io_in_rresp_ready = fringeCommon_io_dram_2_rresp_ready;
  assign MAGToAXI4Bridge_2_io_in_wresp_ready = fringeCommon_io_dram_2_wresp_ready;
  assign MAGToAXI4Bridge_2_io_M_AXI_AWREADY = io_M_AXI_2_AWREADY;
  assign MAGToAXI4Bridge_2_io_M_AXI_ARREADY = io_M_AXI_2_ARREADY;
  assign MAGToAXI4Bridge_2_io_M_AXI_WREADY = io_M_AXI_2_WREADY;
  assign MAGToAXI4Bridge_2_io_M_AXI_RID = io_M_AXI_2_RID;
  assign MAGToAXI4Bridge_2_io_M_AXI_RDATA = io_M_AXI_2_RDATA;
  assign MAGToAXI4Bridge_2_io_M_AXI_RVALID = io_M_AXI_2_RVALID;
  assign MAGToAXI4Bridge_2_io_M_AXI_BID = io_M_AXI_2_BID;
  assign MAGToAXI4Bridge_2_io_M_AXI_BVALID = io_M_AXI_2_BVALID;
  assign MAGToAXI4Bridge_3_io_in_cmd_valid = fringeCommon_io_dram_3_cmd_valid;
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_addr = fringeCommon_io_dram_3_cmd_bits_addr;
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_size = fringeCommon_io_dram_3_cmd_bits_size;
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_isWr = fringeCommon_io_dram_3_cmd_bits_isWr;
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_tag_uid = fringeCommon_io_dram_3_cmd_bits_tag_uid;
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_tag_streamId = fringeCommon_io_dram_3_cmd_bits_tag_streamId;
  assign MAGToAXI4Bridge_3_io_in_wdata_valid = fringeCommon_io_dram_3_wdata_valid;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_3_wdata_bits_wdata_0;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_3_wdata_bits_wdata_1;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_3_wdata_bits_wdata_2;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_3_wdata_bits_wdata_3;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_3_wdata_bits_wdata_4;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_3_wdata_bits_wdata_5;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_3_wdata_bits_wdata_6;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_3_wdata_bits_wdata_7;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_3_wdata_bits_wdata_8;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_3_wdata_bits_wdata_9;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_3_wdata_bits_wdata_10;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_3_wdata_bits_wdata_11;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_3_wdata_bits_wdata_12;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_3_wdata_bits_wdata_13;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_3_wdata_bits_wdata_14;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_3_wdata_bits_wdata_15;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_3_wdata_bits_wstrb_0;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_3_wdata_bits_wstrb_1;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_3_wdata_bits_wstrb_2;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_3_wdata_bits_wstrb_3;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_3_wdata_bits_wstrb_4;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_3_wdata_bits_wstrb_5;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_3_wdata_bits_wstrb_6;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_3_wdata_bits_wstrb_7;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_3_wdata_bits_wstrb_8;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_3_wdata_bits_wstrb_9;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_3_wdata_bits_wstrb_10;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_3_wdata_bits_wstrb_11;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_3_wdata_bits_wstrb_12;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_3_wdata_bits_wstrb_13;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_3_wdata_bits_wstrb_14;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_3_wdata_bits_wstrb_15;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_3_wdata_bits_wstrb_16;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_3_wdata_bits_wstrb_17;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_3_wdata_bits_wstrb_18;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_3_wdata_bits_wstrb_19;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_3_wdata_bits_wstrb_20;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_3_wdata_bits_wstrb_21;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_3_wdata_bits_wstrb_22;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_3_wdata_bits_wstrb_23;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_3_wdata_bits_wstrb_24;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_3_wdata_bits_wstrb_25;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_3_wdata_bits_wstrb_26;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_3_wdata_bits_wstrb_27;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_3_wdata_bits_wstrb_28;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_3_wdata_bits_wstrb_29;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_3_wdata_bits_wstrb_30;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_3_wdata_bits_wstrb_31;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_3_wdata_bits_wstrb_32;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_3_wdata_bits_wstrb_33;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_3_wdata_bits_wstrb_34;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_3_wdata_bits_wstrb_35;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_3_wdata_bits_wstrb_36;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_3_wdata_bits_wstrb_37;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_3_wdata_bits_wstrb_38;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_3_wdata_bits_wstrb_39;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_3_wdata_bits_wstrb_40;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_3_wdata_bits_wstrb_41;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_3_wdata_bits_wstrb_42;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_3_wdata_bits_wstrb_43;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_3_wdata_bits_wstrb_44;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_3_wdata_bits_wstrb_45;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_3_wdata_bits_wstrb_46;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_3_wdata_bits_wstrb_47;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_3_wdata_bits_wstrb_48;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_3_wdata_bits_wstrb_49;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_3_wdata_bits_wstrb_50;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_3_wdata_bits_wstrb_51;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_3_wdata_bits_wstrb_52;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_3_wdata_bits_wstrb_53;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_3_wdata_bits_wstrb_54;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_3_wdata_bits_wstrb_55;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_3_wdata_bits_wstrb_56;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_3_wdata_bits_wstrb_57;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_3_wdata_bits_wstrb_58;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_3_wdata_bits_wstrb_59;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_3_wdata_bits_wstrb_60;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_3_wdata_bits_wstrb_61;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_3_wdata_bits_wstrb_62;
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_3_wdata_bits_wstrb_63;
  assign MAGToAXI4Bridge_3_io_in_rresp_ready = fringeCommon_io_dram_3_rresp_ready;
  assign MAGToAXI4Bridge_3_io_in_wresp_ready = fringeCommon_io_dram_3_wresp_ready;
  assign MAGToAXI4Bridge_3_io_M_AXI_AWREADY = io_M_AXI_3_AWREADY;
  assign MAGToAXI4Bridge_3_io_M_AXI_ARREADY = io_M_AXI_3_ARREADY;
  assign MAGToAXI4Bridge_3_io_M_AXI_WREADY = io_M_AXI_3_WREADY;
  assign MAGToAXI4Bridge_3_io_M_AXI_RID = io_M_AXI_3_RID;
  assign MAGToAXI4Bridge_3_io_M_AXI_RDATA = io_M_AXI_3_RDATA;
  assign MAGToAXI4Bridge_3_io_M_AXI_RVALID = io_M_AXI_3_RVALID;
  assign MAGToAXI4Bridge_3_io_M_AXI_BID = io_M_AXI_3_BID;
  assign MAGToAXI4Bridge_3_io_M_AXI_BVALID = io_M_AXI_3_BVALID;
endmodule
module Top(
  input          clock,
  input          reset,
  input          io_raddr,
  input          io_wen,
  input          io_waddr,
  input          io_wdata,
  output         io_rdata,
  output         io_is_enabled,
  input  [31:0]  io_S_AXI_AWADDR,
  input  [2:0]   io_S_AXI_AWPROT,
  input          io_S_AXI_AWVALID,
  output         io_S_AXI_AWREADY,
  input  [31:0]  io_S_AXI_ARADDR,
  input  [2:0]   io_S_AXI_ARPROT,
  input          io_S_AXI_ARVALID,
  output         io_S_AXI_ARREADY,
  input  [31:0]  io_S_AXI_WDATA,
  input  [3:0]   io_S_AXI_WSTRB,
  input          io_S_AXI_WVALID,
  output         io_S_AXI_WREADY,
  output [31:0]  io_S_AXI_RDATA,
  output [1:0]   io_S_AXI_RRESP,
  output         io_S_AXI_RVALID,
  input          io_S_AXI_RREADY,
  output [1:0]   io_S_AXI_BRESP,
  output         io_S_AXI_BVALID,
  input          io_S_AXI_BREADY,
  output [31:0]  io_M_AXI_0_AWID,
  output [31:0]  io_M_AXI_0_AWUSER,
  output [31:0]  io_M_AXI_0_AWADDR,
  output [7:0]   io_M_AXI_0_AWLEN,
  output [2:0]   io_M_AXI_0_AWSIZE,
  output [1:0]   io_M_AXI_0_AWBURST,
  output         io_M_AXI_0_AWLOCK,
  output [3:0]   io_M_AXI_0_AWCACHE,
  output [2:0]   io_M_AXI_0_AWPROT,
  output [3:0]   io_M_AXI_0_AWQOS,
  output         io_M_AXI_0_AWVALID,
  input          io_M_AXI_0_AWREADY,
  output [31:0]  io_M_AXI_0_ARID,
  output [31:0]  io_M_AXI_0_ARUSER,
  output [31:0]  io_M_AXI_0_ARADDR,
  output [7:0]   io_M_AXI_0_ARLEN,
  output [2:0]   io_M_AXI_0_ARSIZE,
  output [1:0]   io_M_AXI_0_ARBURST,
  output         io_M_AXI_0_ARLOCK,
  output [3:0]   io_M_AXI_0_ARCACHE,
  output [2:0]   io_M_AXI_0_ARPROT,
  output [3:0]   io_M_AXI_0_ARQOS,
  output         io_M_AXI_0_ARVALID,
  input          io_M_AXI_0_ARREADY,
  output [511:0] io_M_AXI_0_WDATA,
  output [63:0]  io_M_AXI_0_WSTRB,
  output         io_M_AXI_0_WLAST,
  output         io_M_AXI_0_WVALID,
  input          io_M_AXI_0_WREADY,
  input  [31:0]  io_M_AXI_0_RID,
  input  [31:0]  io_M_AXI_0_RUSER,
  input  [511:0] io_M_AXI_0_RDATA,
  input  [1:0]   io_M_AXI_0_RRESP,
  input          io_M_AXI_0_RLAST,
  input          io_M_AXI_0_RVALID,
  output         io_M_AXI_0_RREADY,
  input  [31:0]  io_M_AXI_0_BID,
  input  [31:0]  io_M_AXI_0_BUSER,
  input  [1:0]   io_M_AXI_0_BRESP,
  input          io_M_AXI_0_BVALID,
  output         io_M_AXI_0_BREADY,
  output [31:0]  io_M_AXI_1_AWID,
  output [31:0]  io_M_AXI_1_AWUSER,
  output [31:0]  io_M_AXI_1_AWADDR,
  output [7:0]   io_M_AXI_1_AWLEN,
  output [2:0]   io_M_AXI_1_AWSIZE,
  output [1:0]   io_M_AXI_1_AWBURST,
  output         io_M_AXI_1_AWLOCK,
  output [3:0]   io_M_AXI_1_AWCACHE,
  output [2:0]   io_M_AXI_1_AWPROT,
  output [3:0]   io_M_AXI_1_AWQOS,
  output         io_M_AXI_1_AWVALID,
  input          io_M_AXI_1_AWREADY,
  output [31:0]  io_M_AXI_1_ARID,
  output [31:0]  io_M_AXI_1_ARUSER,
  output [31:0]  io_M_AXI_1_ARADDR,
  output [7:0]   io_M_AXI_1_ARLEN,
  output [2:0]   io_M_AXI_1_ARSIZE,
  output [1:0]   io_M_AXI_1_ARBURST,
  output         io_M_AXI_1_ARLOCK,
  output [3:0]   io_M_AXI_1_ARCACHE,
  output [2:0]   io_M_AXI_1_ARPROT,
  output [3:0]   io_M_AXI_1_ARQOS,
  output         io_M_AXI_1_ARVALID,
  input          io_M_AXI_1_ARREADY,
  output [511:0] io_M_AXI_1_WDATA,
  output [63:0]  io_M_AXI_1_WSTRB,
  output         io_M_AXI_1_WLAST,
  output         io_M_AXI_1_WVALID,
  input          io_M_AXI_1_WREADY,
  input  [31:0]  io_M_AXI_1_RID,
  input  [31:0]  io_M_AXI_1_RUSER,
  input  [511:0] io_M_AXI_1_RDATA,
  input  [1:0]   io_M_AXI_1_RRESP,
  input          io_M_AXI_1_RLAST,
  input          io_M_AXI_1_RVALID,
  output         io_M_AXI_1_RREADY,
  input  [31:0]  io_M_AXI_1_BID,
  input  [31:0]  io_M_AXI_1_BUSER,
  input  [1:0]   io_M_AXI_1_BRESP,
  input          io_M_AXI_1_BVALID,
  output         io_M_AXI_1_BREADY,
  output [31:0]  io_M_AXI_2_AWID,
  output [31:0]  io_M_AXI_2_AWUSER,
  output [31:0]  io_M_AXI_2_AWADDR,
  output [7:0]   io_M_AXI_2_AWLEN,
  output [2:0]   io_M_AXI_2_AWSIZE,
  output [1:0]   io_M_AXI_2_AWBURST,
  output         io_M_AXI_2_AWLOCK,
  output [3:0]   io_M_AXI_2_AWCACHE,
  output [2:0]   io_M_AXI_2_AWPROT,
  output [3:0]   io_M_AXI_2_AWQOS,
  output         io_M_AXI_2_AWVALID,
  input          io_M_AXI_2_AWREADY,
  output [31:0]  io_M_AXI_2_ARID,
  output [31:0]  io_M_AXI_2_ARUSER,
  output [31:0]  io_M_AXI_2_ARADDR,
  output [7:0]   io_M_AXI_2_ARLEN,
  output [2:0]   io_M_AXI_2_ARSIZE,
  output [1:0]   io_M_AXI_2_ARBURST,
  output         io_M_AXI_2_ARLOCK,
  output [3:0]   io_M_AXI_2_ARCACHE,
  output [2:0]   io_M_AXI_2_ARPROT,
  output [3:0]   io_M_AXI_2_ARQOS,
  output         io_M_AXI_2_ARVALID,
  input          io_M_AXI_2_ARREADY,
  output [511:0] io_M_AXI_2_WDATA,
  output [63:0]  io_M_AXI_2_WSTRB,
  output         io_M_AXI_2_WLAST,
  output         io_M_AXI_2_WVALID,
  input          io_M_AXI_2_WREADY,
  input  [31:0]  io_M_AXI_2_RID,
  input  [31:0]  io_M_AXI_2_RUSER,
  input  [511:0] io_M_AXI_2_RDATA,
  input  [1:0]   io_M_AXI_2_RRESP,
  input          io_M_AXI_2_RLAST,
  input          io_M_AXI_2_RVALID,
  output         io_M_AXI_2_RREADY,
  input  [31:0]  io_M_AXI_2_BID,
  input  [31:0]  io_M_AXI_2_BUSER,
  input  [1:0]   io_M_AXI_2_BRESP,
  input          io_M_AXI_2_BVALID,
  output         io_M_AXI_2_BREADY,
  output [31:0]  io_M_AXI_3_AWID,
  output [31:0]  io_M_AXI_3_AWUSER,
  output [31:0]  io_M_AXI_3_AWADDR,
  output [7:0]   io_M_AXI_3_AWLEN,
  output [2:0]   io_M_AXI_3_AWSIZE,
  output [1:0]   io_M_AXI_3_AWBURST,
  output         io_M_AXI_3_AWLOCK,
  output [3:0]   io_M_AXI_3_AWCACHE,
  output [2:0]   io_M_AXI_3_AWPROT,
  output [3:0]   io_M_AXI_3_AWQOS,
  output         io_M_AXI_3_AWVALID,
  input          io_M_AXI_3_AWREADY,
  output [31:0]  io_M_AXI_3_ARID,
  output [31:0]  io_M_AXI_3_ARUSER,
  output [31:0]  io_M_AXI_3_ARADDR,
  output [7:0]   io_M_AXI_3_ARLEN,
  output [2:0]   io_M_AXI_3_ARSIZE,
  output [1:0]   io_M_AXI_3_ARBURST,
  output         io_M_AXI_3_ARLOCK,
  output [3:0]   io_M_AXI_3_ARCACHE,
  output [2:0]   io_M_AXI_3_ARPROT,
  output [3:0]   io_M_AXI_3_ARQOS,
  output         io_M_AXI_3_ARVALID,
  input          io_M_AXI_3_ARREADY,
  output [511:0] io_M_AXI_3_WDATA,
  output [63:0]  io_M_AXI_3_WSTRB,
  output         io_M_AXI_3_WLAST,
  output         io_M_AXI_3_WVALID,
  input          io_M_AXI_3_WREADY,
  input  [31:0]  io_M_AXI_3_RID,
  input  [31:0]  io_M_AXI_3_RUSER,
  input  [511:0] io_M_AXI_3_RDATA,
  input  [1:0]   io_M_AXI_3_RRESP,
  input          io_M_AXI_3_RLAST,
  input          io_M_AXI_3_RVALID,
  output         io_M_AXI_3_RREADY,
  input  [31:0]  io_M_AXI_3_BID,
  input  [31:0]  io_M_AXI_3_BUSER,
  input  [1:0]   io_M_AXI_3_BRESP,
  input          io_M_AXI_3_BVALID,
  output         io_M_AXI_3_BREADY,
  input          io_TOP_AXI_AWID,
  input  [31:0]  io_TOP_AXI_AWUSER,
  input  [31:0]  io_TOP_AXI_AWADDR,
  input  [7:0]   io_TOP_AXI_AWLEN,
  input  [2:0]   io_TOP_AXI_AWSIZE,
  input  [1:0]   io_TOP_AXI_AWBURST,
  input          io_TOP_AXI_AWLOCK,
  input  [3:0]   io_TOP_AXI_AWCACHE,
  input  [2:0]   io_TOP_AXI_AWPROT,
  input  [3:0]   io_TOP_AXI_AWQOS,
  input          io_TOP_AXI_AWVALID,
  input          io_TOP_AXI_AWREADY,
  input          io_TOP_AXI_ARID,
  input  [31:0]  io_TOP_AXI_ARUSER,
  input  [31:0]  io_TOP_AXI_ARADDR,
  input  [7:0]   io_TOP_AXI_ARLEN,
  input  [2:0]   io_TOP_AXI_ARSIZE,
  input  [1:0]   io_TOP_AXI_ARBURST,
  input          io_TOP_AXI_ARLOCK,
  input  [3:0]   io_TOP_AXI_ARCACHE,
  input  [2:0]   io_TOP_AXI_ARPROT,
  input  [3:0]   io_TOP_AXI_ARQOS,
  input          io_TOP_AXI_ARVALID,
  input          io_TOP_AXI_ARREADY,
  input  [31:0]  io_TOP_AXI_WDATA,
  input  [63:0]  io_TOP_AXI_WSTRB,
  input          io_TOP_AXI_WLAST,
  input          io_TOP_AXI_WVALID,
  input          io_TOP_AXI_WREADY,
  input          io_TOP_AXI_RID,
  input  [31:0]  io_TOP_AXI_RUSER,
  input  [31:0]  io_TOP_AXI_RDATA,
  input  [1:0]   io_TOP_AXI_RRESP,
  input          io_TOP_AXI_RLAST,
  input          io_TOP_AXI_RVALID,
  input          io_TOP_AXI_RREADY,
  input          io_TOP_AXI_BID,
  input  [31:0]  io_TOP_AXI_BUSER,
  input  [1:0]   io_TOP_AXI_BRESP,
  input          io_TOP_AXI_BVALID,
  input          io_TOP_AXI_BREADY,
  input          io_DWIDTH_AXI_AWID,
  input  [31:0]  io_DWIDTH_AXI_AWUSER,
  input  [31:0]  io_DWIDTH_AXI_AWADDR,
  input  [7:0]   io_DWIDTH_AXI_AWLEN,
  input  [2:0]   io_DWIDTH_AXI_AWSIZE,
  input  [1:0]   io_DWIDTH_AXI_AWBURST,
  input          io_DWIDTH_AXI_AWLOCK,
  input  [3:0]   io_DWIDTH_AXI_AWCACHE,
  input  [2:0]   io_DWIDTH_AXI_AWPROT,
  input  [3:0]   io_DWIDTH_AXI_AWQOS,
  input          io_DWIDTH_AXI_AWVALID,
  input          io_DWIDTH_AXI_AWREADY,
  input          io_DWIDTH_AXI_ARID,
  input  [31:0]  io_DWIDTH_AXI_ARUSER,
  input  [31:0]  io_DWIDTH_AXI_ARADDR,
  input  [7:0]   io_DWIDTH_AXI_ARLEN,
  input  [2:0]   io_DWIDTH_AXI_ARSIZE,
  input  [1:0]   io_DWIDTH_AXI_ARBURST,
  input          io_DWIDTH_AXI_ARLOCK,
  input  [3:0]   io_DWIDTH_AXI_ARCACHE,
  input  [2:0]   io_DWIDTH_AXI_ARPROT,
  input  [3:0]   io_DWIDTH_AXI_ARQOS,
  input          io_DWIDTH_AXI_ARVALID,
  input          io_DWIDTH_AXI_ARREADY,
  input  [31:0]  io_DWIDTH_AXI_WDATA,
  input  [63:0]  io_DWIDTH_AXI_WSTRB,
  input          io_DWIDTH_AXI_WLAST,
  input          io_DWIDTH_AXI_WVALID,
  input          io_DWIDTH_AXI_WREADY,
  input          io_DWIDTH_AXI_RID,
  input  [31:0]  io_DWIDTH_AXI_RUSER,
  input  [31:0]  io_DWIDTH_AXI_RDATA,
  input  [1:0]   io_DWIDTH_AXI_RRESP,
  input          io_DWIDTH_AXI_RLAST,
  input          io_DWIDTH_AXI_RVALID,
  input          io_DWIDTH_AXI_RREADY,
  input          io_DWIDTH_AXI_BID,
  input  [31:0]  io_DWIDTH_AXI_BUSER,
  input  [1:0]   io_DWIDTH_AXI_BRESP,
  input          io_DWIDTH_AXI_BVALID,
  input          io_DWIDTH_AXI_BREADY,
  input          io_PROTOCOL_AXI_AWID,
  input  [31:0]  io_PROTOCOL_AXI_AWUSER,
  input  [31:0]  io_PROTOCOL_AXI_AWADDR,
  input  [7:0]   io_PROTOCOL_AXI_AWLEN,
  input  [2:0]   io_PROTOCOL_AXI_AWSIZE,
  input  [1:0]   io_PROTOCOL_AXI_AWBURST,
  input          io_PROTOCOL_AXI_AWLOCK,
  input  [3:0]   io_PROTOCOL_AXI_AWCACHE,
  input  [2:0]   io_PROTOCOL_AXI_AWPROT,
  input  [3:0]   io_PROTOCOL_AXI_AWQOS,
  input          io_PROTOCOL_AXI_AWVALID,
  input          io_PROTOCOL_AXI_AWREADY,
  input          io_PROTOCOL_AXI_ARID,
  input  [31:0]  io_PROTOCOL_AXI_ARUSER,
  input  [31:0]  io_PROTOCOL_AXI_ARADDR,
  input  [7:0]   io_PROTOCOL_AXI_ARLEN,
  input  [2:0]   io_PROTOCOL_AXI_ARSIZE,
  input  [1:0]   io_PROTOCOL_AXI_ARBURST,
  input          io_PROTOCOL_AXI_ARLOCK,
  input  [3:0]   io_PROTOCOL_AXI_ARCACHE,
  input  [2:0]   io_PROTOCOL_AXI_ARPROT,
  input  [3:0]   io_PROTOCOL_AXI_ARQOS,
  input          io_PROTOCOL_AXI_ARVALID,
  input          io_PROTOCOL_AXI_ARREADY,
  input  [31:0]  io_PROTOCOL_AXI_WDATA,
  input  [63:0]  io_PROTOCOL_AXI_WSTRB,
  input          io_PROTOCOL_AXI_WLAST,
  input          io_PROTOCOL_AXI_WVALID,
  input          io_PROTOCOL_AXI_WREADY,
  input          io_PROTOCOL_AXI_RID,
  input  [31:0]  io_PROTOCOL_AXI_RUSER,
  input  [31:0]  io_PROTOCOL_AXI_RDATA,
  input  [1:0]   io_PROTOCOL_AXI_RRESP,
  input          io_PROTOCOL_AXI_RLAST,
  input          io_PROTOCOL_AXI_RVALID,
  input          io_PROTOCOL_AXI_RREADY,
  input          io_PROTOCOL_AXI_BID,
  input  [31:0]  io_PROTOCOL_AXI_BUSER,
  input  [1:0]   io_PROTOCOL_AXI_BRESP,
  input          io_PROTOCOL_AXI_BVALID,
  input          io_PROTOCOL_AXI_BREADY,
  input          io_CLOCKCONVERT_AXI_AWID,
  input  [31:0]  io_CLOCKCONVERT_AXI_AWUSER,
  input  [31:0]  io_CLOCKCONVERT_AXI_AWADDR,
  input  [7:0]   io_CLOCKCONVERT_AXI_AWLEN,
  input  [2:0]   io_CLOCKCONVERT_AXI_AWSIZE,
  input  [1:0]   io_CLOCKCONVERT_AXI_AWBURST,
  input          io_CLOCKCONVERT_AXI_AWLOCK,
  input  [3:0]   io_CLOCKCONVERT_AXI_AWCACHE,
  input  [2:0]   io_CLOCKCONVERT_AXI_AWPROT,
  input  [3:0]   io_CLOCKCONVERT_AXI_AWQOS,
  input          io_CLOCKCONVERT_AXI_AWVALID,
  input          io_CLOCKCONVERT_AXI_AWREADY,
  input          io_CLOCKCONVERT_AXI_ARID,
  input  [31:0]  io_CLOCKCONVERT_AXI_ARUSER,
  input  [31:0]  io_CLOCKCONVERT_AXI_ARADDR,
  input  [7:0]   io_CLOCKCONVERT_AXI_ARLEN,
  input  [2:0]   io_CLOCKCONVERT_AXI_ARSIZE,
  input  [1:0]   io_CLOCKCONVERT_AXI_ARBURST,
  input          io_CLOCKCONVERT_AXI_ARLOCK,
  input  [3:0]   io_CLOCKCONVERT_AXI_ARCACHE,
  input  [2:0]   io_CLOCKCONVERT_AXI_ARPROT,
  input  [3:0]   io_CLOCKCONVERT_AXI_ARQOS,
  input          io_CLOCKCONVERT_AXI_ARVALID,
  input          io_CLOCKCONVERT_AXI_ARREADY,
  input  [31:0]  io_CLOCKCONVERT_AXI_WDATA,
  input  [63:0]  io_CLOCKCONVERT_AXI_WSTRB,
  input          io_CLOCKCONVERT_AXI_WLAST,
  input          io_CLOCKCONVERT_AXI_WVALID,
  input          io_CLOCKCONVERT_AXI_WREADY,
  input          io_CLOCKCONVERT_AXI_RID,
  input  [31:0]  io_CLOCKCONVERT_AXI_RUSER,
  input  [31:0]  io_CLOCKCONVERT_AXI_RDATA,
  input  [1:0]   io_CLOCKCONVERT_AXI_RRESP,
  input          io_CLOCKCONVERT_AXI_RLAST,
  input          io_CLOCKCONVERT_AXI_RVALID,
  input          io_CLOCKCONVERT_AXI_RREADY,
  input          io_CLOCKCONVERT_AXI_BID,
  input  [31:0]  io_CLOCKCONVERT_AXI_BUSER,
  input  [1:0]   io_CLOCKCONVERT_AXI_BRESP,
  input          io_CLOCKCONVERT_AXI_BVALID,
  input          io_CLOCKCONVERT_AXI_BREADY
);
  wire  accel_clock;
  wire  accel_reset;
  wire  accel_io_enable;
  wire  accel_io_done;
  wire  accel_io_memStreams_loads_3_cmd_ready;
  wire  accel_io_memStreams_loads_3_cmd_valid;
  wire [63:0] accel_io_memStreams_loads_3_cmd_bits_addr;
  wire  accel_io_memStreams_loads_3_cmd_bits_isWr;
  wire [15:0] accel_io_memStreams_loads_3_cmd_bits_size;
  wire  accel_io_memStreams_loads_3_rdata_ready;
  wire  accel_io_memStreams_loads_3_rdata_valid;
  wire [31:0] accel_io_memStreams_loads_3_rdata_bits_0;
  wire  accel_io_memStreams_loads_2_cmd_ready;
  wire  accel_io_memStreams_loads_2_cmd_valid;
  wire [63:0] accel_io_memStreams_loads_2_cmd_bits_addr;
  wire  accel_io_memStreams_loads_2_cmd_bits_isWr;
  wire [15:0] accel_io_memStreams_loads_2_cmd_bits_size;
  wire  accel_io_memStreams_loads_2_rdata_ready;
  wire  accel_io_memStreams_loads_2_rdata_valid;
  wire [31:0] accel_io_memStreams_loads_2_rdata_bits_0;
  wire  accel_io_memStreams_loads_1_cmd_ready;
  wire  accel_io_memStreams_loads_1_cmd_valid;
  wire [63:0] accel_io_memStreams_loads_1_cmd_bits_addr;
  wire  accel_io_memStreams_loads_1_cmd_bits_isWr;
  wire [15:0] accel_io_memStreams_loads_1_cmd_bits_size;
  wire  accel_io_memStreams_loads_1_rdata_ready;
  wire  accel_io_memStreams_loads_1_rdata_valid;
  wire [31:0] accel_io_memStreams_loads_1_rdata_bits_0;
  wire  accel_io_memStreams_loads_0_cmd_ready;
  wire  accel_io_memStreams_loads_0_cmd_valid;
  wire [63:0] accel_io_memStreams_loads_0_cmd_bits_addr;
  wire  accel_io_memStreams_loads_0_cmd_bits_isWr;
  wire [15:0] accel_io_memStreams_loads_0_cmd_bits_size;
  wire  accel_io_memStreams_loads_0_rdata_ready;
  wire  accel_io_memStreams_loads_0_rdata_valid;
  wire [31:0] accel_io_memStreams_loads_0_rdata_bits_0;
  wire [63:0] accel_io_argIns_0;
  wire [63:0] accel_io_argIns_1;
  wire [63:0] accel_io_argIns_2;
  wire  accel_io_argOuts_0_valid;
  wire [63:0] accel_io_argOuts_0_bits;
  wire  FringeZynq_clock;
  wire  FringeZynq_reset;
  wire [31:0] FringeZynq_io_S_AXI_AWADDR;
  wire [2:0] FringeZynq_io_S_AXI_AWPROT;
  wire  FringeZynq_io_S_AXI_AWVALID;
  wire  FringeZynq_io_S_AXI_AWREADY;
  wire [31:0] FringeZynq_io_S_AXI_ARADDR;
  wire [2:0] FringeZynq_io_S_AXI_ARPROT;
  wire  FringeZynq_io_S_AXI_ARVALID;
  wire  FringeZynq_io_S_AXI_ARREADY;
  wire [31:0] FringeZynq_io_S_AXI_WDATA;
  wire [3:0] FringeZynq_io_S_AXI_WSTRB;
  wire  FringeZynq_io_S_AXI_WVALID;
  wire  FringeZynq_io_S_AXI_WREADY;
  wire [31:0] FringeZynq_io_S_AXI_RDATA;
  wire [1:0] FringeZynq_io_S_AXI_RRESP;
  wire  FringeZynq_io_S_AXI_RVALID;
  wire  FringeZynq_io_S_AXI_RREADY;
  wire [1:0] FringeZynq_io_S_AXI_BRESP;
  wire  FringeZynq_io_S_AXI_BVALID;
  wire  FringeZynq_io_S_AXI_BREADY;
  wire [31:0] FringeZynq_io_M_AXI_0_AWID;
  wire [31:0] FringeZynq_io_M_AXI_0_AWADDR;
  wire [7:0] FringeZynq_io_M_AXI_0_AWLEN;
  wire  FringeZynq_io_M_AXI_0_AWVALID;
  wire  FringeZynq_io_M_AXI_0_AWREADY;
  wire [31:0] FringeZynq_io_M_AXI_0_ARID;
  wire [31:0] FringeZynq_io_M_AXI_0_ARADDR;
  wire [7:0] FringeZynq_io_M_AXI_0_ARLEN;
  wire  FringeZynq_io_M_AXI_0_ARVALID;
  wire  FringeZynq_io_M_AXI_0_ARREADY;
  wire [511:0] FringeZynq_io_M_AXI_0_WDATA;
  wire [63:0] FringeZynq_io_M_AXI_0_WSTRB;
  wire  FringeZynq_io_M_AXI_0_WVALID;
  wire  FringeZynq_io_M_AXI_0_WREADY;
  wire [31:0] FringeZynq_io_M_AXI_0_RID;
  wire [511:0] FringeZynq_io_M_AXI_0_RDATA;
  wire  FringeZynq_io_M_AXI_0_RVALID;
  wire  FringeZynq_io_M_AXI_0_RREADY;
  wire [31:0] FringeZynq_io_M_AXI_0_BID;
  wire  FringeZynq_io_M_AXI_0_BVALID;
  wire  FringeZynq_io_M_AXI_0_BREADY;
  wire [31:0] FringeZynq_io_M_AXI_1_AWID;
  wire [31:0] FringeZynq_io_M_AXI_1_AWADDR;
  wire [7:0] FringeZynq_io_M_AXI_1_AWLEN;
  wire  FringeZynq_io_M_AXI_1_AWVALID;
  wire  FringeZynq_io_M_AXI_1_AWREADY;
  wire [31:0] FringeZynq_io_M_AXI_1_ARID;
  wire [31:0] FringeZynq_io_M_AXI_1_ARADDR;
  wire [7:0] FringeZynq_io_M_AXI_1_ARLEN;
  wire  FringeZynq_io_M_AXI_1_ARVALID;
  wire  FringeZynq_io_M_AXI_1_ARREADY;
  wire [511:0] FringeZynq_io_M_AXI_1_WDATA;
  wire [63:0] FringeZynq_io_M_AXI_1_WSTRB;
  wire  FringeZynq_io_M_AXI_1_WVALID;
  wire  FringeZynq_io_M_AXI_1_WREADY;
  wire [31:0] FringeZynq_io_M_AXI_1_RID;
  wire [511:0] FringeZynq_io_M_AXI_1_RDATA;
  wire  FringeZynq_io_M_AXI_1_RVALID;
  wire  FringeZynq_io_M_AXI_1_RREADY;
  wire [31:0] FringeZynq_io_M_AXI_1_BID;
  wire  FringeZynq_io_M_AXI_1_BVALID;
  wire  FringeZynq_io_M_AXI_1_BREADY;
  wire [31:0] FringeZynq_io_M_AXI_2_AWID;
  wire [31:0] FringeZynq_io_M_AXI_2_AWADDR;
  wire [7:0] FringeZynq_io_M_AXI_2_AWLEN;
  wire  FringeZynq_io_M_AXI_2_AWVALID;
  wire  FringeZynq_io_M_AXI_2_AWREADY;
  wire [31:0] FringeZynq_io_M_AXI_2_ARID;
  wire [31:0] FringeZynq_io_M_AXI_2_ARADDR;
  wire [7:0] FringeZynq_io_M_AXI_2_ARLEN;
  wire  FringeZynq_io_M_AXI_2_ARVALID;
  wire  FringeZynq_io_M_AXI_2_ARREADY;
  wire [511:0] FringeZynq_io_M_AXI_2_WDATA;
  wire [63:0] FringeZynq_io_M_AXI_2_WSTRB;
  wire  FringeZynq_io_M_AXI_2_WVALID;
  wire  FringeZynq_io_M_AXI_2_WREADY;
  wire [31:0] FringeZynq_io_M_AXI_2_RID;
  wire [511:0] FringeZynq_io_M_AXI_2_RDATA;
  wire  FringeZynq_io_M_AXI_2_RVALID;
  wire  FringeZynq_io_M_AXI_2_RREADY;
  wire [31:0] FringeZynq_io_M_AXI_2_BID;
  wire  FringeZynq_io_M_AXI_2_BVALID;
  wire  FringeZynq_io_M_AXI_2_BREADY;
  wire [31:0] FringeZynq_io_M_AXI_3_AWID;
  wire [31:0] FringeZynq_io_M_AXI_3_AWADDR;
  wire [7:0] FringeZynq_io_M_AXI_3_AWLEN;
  wire  FringeZynq_io_M_AXI_3_AWVALID;
  wire  FringeZynq_io_M_AXI_3_AWREADY;
  wire [31:0] FringeZynq_io_M_AXI_3_ARID;
  wire [31:0] FringeZynq_io_M_AXI_3_ARADDR;
  wire [7:0] FringeZynq_io_M_AXI_3_ARLEN;
  wire  FringeZynq_io_M_AXI_3_ARVALID;
  wire  FringeZynq_io_M_AXI_3_ARREADY;
  wire [511:0] FringeZynq_io_M_AXI_3_WDATA;
  wire [63:0] FringeZynq_io_M_AXI_3_WSTRB;
  wire  FringeZynq_io_M_AXI_3_WVALID;
  wire  FringeZynq_io_M_AXI_3_WREADY;
  wire [31:0] FringeZynq_io_M_AXI_3_RID;
  wire [511:0] FringeZynq_io_M_AXI_3_RDATA;
  wire  FringeZynq_io_M_AXI_3_RVALID;
  wire  FringeZynq_io_M_AXI_3_RREADY;
  wire [31:0] FringeZynq_io_M_AXI_3_BID;
  wire  FringeZynq_io_M_AXI_3_BVALID;
  wire  FringeZynq_io_M_AXI_3_BREADY;
  wire [31:0] FringeZynq_io_TOP_AXI_AWADDR;
  wire [7:0] FringeZynq_io_TOP_AXI_AWLEN;
  wire  FringeZynq_io_TOP_AXI_AWVALID;
  wire  FringeZynq_io_TOP_AXI_AWREADY;
  wire  FringeZynq_io_TOP_AXI_ARID;
  wire [31:0] FringeZynq_io_TOP_AXI_ARADDR;
  wire [7:0] FringeZynq_io_TOP_AXI_ARLEN;
  wire [2:0] FringeZynq_io_TOP_AXI_ARSIZE;
  wire [1:0] FringeZynq_io_TOP_AXI_ARBURST;
  wire  FringeZynq_io_TOP_AXI_ARVALID;
  wire  FringeZynq_io_TOP_AXI_ARREADY;
  wire [31:0] FringeZynq_io_TOP_AXI_WDATA;
  wire [63:0] FringeZynq_io_TOP_AXI_WSTRB;
  wire  FringeZynq_io_TOP_AXI_WVALID;
  wire  FringeZynq_io_TOP_AXI_WREADY;
  wire  FringeZynq_io_TOP_AXI_RVALID;
  wire  FringeZynq_io_TOP_AXI_RREADY;
  wire  FringeZynq_io_TOP_AXI_BVALID;
  wire  FringeZynq_io_TOP_AXI_BREADY;
  wire [31:0] FringeZynq_io_DWIDTH_AXI_AWADDR;
  wire [7:0] FringeZynq_io_DWIDTH_AXI_AWLEN;
  wire  FringeZynq_io_DWIDTH_AXI_AWVALID;
  wire  FringeZynq_io_DWIDTH_AXI_AWREADY;
  wire [31:0] FringeZynq_io_DWIDTH_AXI_ARADDR;
  wire [7:0] FringeZynq_io_DWIDTH_AXI_ARLEN;
  wire [2:0] FringeZynq_io_DWIDTH_AXI_ARSIZE;
  wire [1:0] FringeZynq_io_DWIDTH_AXI_ARBURST;
  wire  FringeZynq_io_DWIDTH_AXI_ARVALID;
  wire  FringeZynq_io_DWIDTH_AXI_ARREADY;
  wire [31:0] FringeZynq_io_DWIDTH_AXI_WDATA;
  wire [63:0] FringeZynq_io_DWIDTH_AXI_WSTRB;
  wire  FringeZynq_io_DWIDTH_AXI_WVALID;
  wire  FringeZynq_io_DWIDTH_AXI_WREADY;
  wire  FringeZynq_io_DWIDTH_AXI_RVALID;
  wire  FringeZynq_io_DWIDTH_AXI_RREADY;
  wire  FringeZynq_io_DWIDTH_AXI_BVALID;
  wire  FringeZynq_io_DWIDTH_AXI_BREADY;
  wire  FringeZynq_io_enable;
  wire  FringeZynq_io_done;
  wire  FringeZynq_io_reset;
  wire [63:0] FringeZynq_io_argIns_0;
  wire [63:0] FringeZynq_io_argIns_1;
  wire [63:0] FringeZynq_io_argIns_2;
  wire  FringeZynq_io_argOuts_0_valid;
  wire [63:0] FringeZynq_io_argOuts_0_bits;
  wire  FringeZynq_io_memStreams_loads_3_cmd_ready;
  wire  FringeZynq_io_memStreams_loads_3_cmd_valid;
  wire [63:0] FringeZynq_io_memStreams_loads_3_cmd_bits_addr;
  wire  FringeZynq_io_memStreams_loads_3_cmd_bits_isWr;
  wire [15:0] FringeZynq_io_memStreams_loads_3_cmd_bits_size;
  wire  FringeZynq_io_memStreams_loads_3_rdata_ready;
  wire  FringeZynq_io_memStreams_loads_3_rdata_valid;
  wire [31:0] FringeZynq_io_memStreams_loads_3_rdata_bits_0;
  wire  FringeZynq_io_memStreams_loads_2_cmd_ready;
  wire  FringeZynq_io_memStreams_loads_2_cmd_valid;
  wire [63:0] FringeZynq_io_memStreams_loads_2_cmd_bits_addr;
  wire  FringeZynq_io_memStreams_loads_2_cmd_bits_isWr;
  wire [15:0] FringeZynq_io_memStreams_loads_2_cmd_bits_size;
  wire  FringeZynq_io_memStreams_loads_2_rdata_ready;
  wire  FringeZynq_io_memStreams_loads_2_rdata_valid;
  wire [31:0] FringeZynq_io_memStreams_loads_2_rdata_bits_0;
  wire  FringeZynq_io_memStreams_loads_1_cmd_ready;
  wire  FringeZynq_io_memStreams_loads_1_cmd_valid;
  wire [63:0] FringeZynq_io_memStreams_loads_1_cmd_bits_addr;
  wire  FringeZynq_io_memStreams_loads_1_cmd_bits_isWr;
  wire [15:0] FringeZynq_io_memStreams_loads_1_cmd_bits_size;
  wire  FringeZynq_io_memStreams_loads_1_rdata_ready;
  wire  FringeZynq_io_memStreams_loads_1_rdata_valid;
  wire [31:0] FringeZynq_io_memStreams_loads_1_rdata_bits_0;
  wire  FringeZynq_io_memStreams_loads_0_cmd_ready;
  wire  FringeZynq_io_memStreams_loads_0_cmd_valid;
  wire [63:0] FringeZynq_io_memStreams_loads_0_cmd_bits_addr;
  wire  FringeZynq_io_memStreams_loads_0_cmd_bits_isWr;
  wire [15:0] FringeZynq_io_memStreams_loads_0_cmd_bits_size;
  wire  FringeZynq_io_memStreams_loads_0_rdata_ready;
  wire  FringeZynq_io_memStreams_loads_0_rdata_valid;
  wire [31:0] FringeZynq_io_memStreams_loads_0_rdata_bits_0;
  wire  _T_475;
  wire  _T_476;
  AccelTop accel (
    .clock(accel_clock),
    .reset(accel_reset),
    .io_enable(accel_io_enable),
    .io_done(accel_io_done),
    .io_memStreams_loads_3_cmd_ready(accel_io_memStreams_loads_3_cmd_ready),
    .io_memStreams_loads_3_cmd_valid(accel_io_memStreams_loads_3_cmd_valid),
    .io_memStreams_loads_3_cmd_bits_addr(accel_io_memStreams_loads_3_cmd_bits_addr),
    .io_memStreams_loads_3_cmd_bits_isWr(accel_io_memStreams_loads_3_cmd_bits_isWr),
    .io_memStreams_loads_3_cmd_bits_size(accel_io_memStreams_loads_3_cmd_bits_size),
    .io_memStreams_loads_3_rdata_ready(accel_io_memStreams_loads_3_rdata_ready),
    .io_memStreams_loads_3_rdata_valid(accel_io_memStreams_loads_3_rdata_valid),
    .io_memStreams_loads_3_rdata_bits_0(accel_io_memStreams_loads_3_rdata_bits_0),
    .io_memStreams_loads_2_cmd_ready(accel_io_memStreams_loads_2_cmd_ready),
    .io_memStreams_loads_2_cmd_valid(accel_io_memStreams_loads_2_cmd_valid),
    .io_memStreams_loads_2_cmd_bits_addr(accel_io_memStreams_loads_2_cmd_bits_addr),
    .io_memStreams_loads_2_cmd_bits_isWr(accel_io_memStreams_loads_2_cmd_bits_isWr),
    .io_memStreams_loads_2_cmd_bits_size(accel_io_memStreams_loads_2_cmd_bits_size),
    .io_memStreams_loads_2_rdata_ready(accel_io_memStreams_loads_2_rdata_ready),
    .io_memStreams_loads_2_rdata_valid(accel_io_memStreams_loads_2_rdata_valid),
    .io_memStreams_loads_2_rdata_bits_0(accel_io_memStreams_loads_2_rdata_bits_0),
    .io_memStreams_loads_1_cmd_ready(accel_io_memStreams_loads_1_cmd_ready),
    .io_memStreams_loads_1_cmd_valid(accel_io_memStreams_loads_1_cmd_valid),
    .io_memStreams_loads_1_cmd_bits_addr(accel_io_memStreams_loads_1_cmd_bits_addr),
    .io_memStreams_loads_1_cmd_bits_isWr(accel_io_memStreams_loads_1_cmd_bits_isWr),
    .io_memStreams_loads_1_cmd_bits_size(accel_io_memStreams_loads_1_cmd_bits_size),
    .io_memStreams_loads_1_rdata_ready(accel_io_memStreams_loads_1_rdata_ready),
    .io_memStreams_loads_1_rdata_valid(accel_io_memStreams_loads_1_rdata_valid),
    .io_memStreams_loads_1_rdata_bits_0(accel_io_memStreams_loads_1_rdata_bits_0),
    .io_memStreams_loads_0_cmd_ready(accel_io_memStreams_loads_0_cmd_ready),
    .io_memStreams_loads_0_cmd_valid(accel_io_memStreams_loads_0_cmd_valid),
    .io_memStreams_loads_0_cmd_bits_addr(accel_io_memStreams_loads_0_cmd_bits_addr),
    .io_memStreams_loads_0_cmd_bits_isWr(accel_io_memStreams_loads_0_cmd_bits_isWr),
    .io_memStreams_loads_0_cmd_bits_size(accel_io_memStreams_loads_0_cmd_bits_size),
    .io_memStreams_loads_0_rdata_ready(accel_io_memStreams_loads_0_rdata_ready),
    .io_memStreams_loads_0_rdata_valid(accel_io_memStreams_loads_0_rdata_valid),
    .io_memStreams_loads_0_rdata_bits_0(accel_io_memStreams_loads_0_rdata_bits_0),
    .io_argIns_0(accel_io_argIns_0),
    .io_argIns_1(accel_io_argIns_1),
    .io_argIns_2(accel_io_argIns_2),
    .io_argOuts_0_valid(accel_io_argOuts_0_valid),
    .io_argOuts_0_bits(accel_io_argOuts_0_bits)
  );
  FringeZynq FringeZynq (
    .clock(FringeZynq_clock),
    .reset(FringeZynq_reset),
    .io_S_AXI_AWADDR(FringeZynq_io_S_AXI_AWADDR),
    .io_S_AXI_AWPROT(FringeZynq_io_S_AXI_AWPROT),
    .io_S_AXI_AWVALID(FringeZynq_io_S_AXI_AWVALID),
    .io_S_AXI_AWREADY(FringeZynq_io_S_AXI_AWREADY),
    .io_S_AXI_ARADDR(FringeZynq_io_S_AXI_ARADDR),
    .io_S_AXI_ARPROT(FringeZynq_io_S_AXI_ARPROT),
    .io_S_AXI_ARVALID(FringeZynq_io_S_AXI_ARVALID),
    .io_S_AXI_ARREADY(FringeZynq_io_S_AXI_ARREADY),
    .io_S_AXI_WDATA(FringeZynq_io_S_AXI_WDATA),
    .io_S_AXI_WSTRB(FringeZynq_io_S_AXI_WSTRB),
    .io_S_AXI_WVALID(FringeZynq_io_S_AXI_WVALID),
    .io_S_AXI_WREADY(FringeZynq_io_S_AXI_WREADY),
    .io_S_AXI_RDATA(FringeZynq_io_S_AXI_RDATA),
    .io_S_AXI_RRESP(FringeZynq_io_S_AXI_RRESP),
    .io_S_AXI_RVALID(FringeZynq_io_S_AXI_RVALID),
    .io_S_AXI_RREADY(FringeZynq_io_S_AXI_RREADY),
    .io_S_AXI_BRESP(FringeZynq_io_S_AXI_BRESP),
    .io_S_AXI_BVALID(FringeZynq_io_S_AXI_BVALID),
    .io_S_AXI_BREADY(FringeZynq_io_S_AXI_BREADY),
    .io_M_AXI_0_AWID(FringeZynq_io_M_AXI_0_AWID),
    .io_M_AXI_0_AWADDR(FringeZynq_io_M_AXI_0_AWADDR),
    .io_M_AXI_0_AWLEN(FringeZynq_io_M_AXI_0_AWLEN),
    .io_M_AXI_0_AWVALID(FringeZynq_io_M_AXI_0_AWVALID),
    .io_M_AXI_0_AWREADY(FringeZynq_io_M_AXI_0_AWREADY),
    .io_M_AXI_0_ARID(FringeZynq_io_M_AXI_0_ARID),
    .io_M_AXI_0_ARADDR(FringeZynq_io_M_AXI_0_ARADDR),
    .io_M_AXI_0_ARLEN(FringeZynq_io_M_AXI_0_ARLEN),
    .io_M_AXI_0_ARVALID(FringeZynq_io_M_AXI_0_ARVALID),
    .io_M_AXI_0_ARREADY(FringeZynq_io_M_AXI_0_ARREADY),
    .io_M_AXI_0_WDATA(FringeZynq_io_M_AXI_0_WDATA),
    .io_M_AXI_0_WSTRB(FringeZynq_io_M_AXI_0_WSTRB),
    .io_M_AXI_0_WVALID(FringeZynq_io_M_AXI_0_WVALID),
    .io_M_AXI_0_WREADY(FringeZynq_io_M_AXI_0_WREADY),
    .io_M_AXI_0_RID(FringeZynq_io_M_AXI_0_RID),
    .io_M_AXI_0_RDATA(FringeZynq_io_M_AXI_0_RDATA),
    .io_M_AXI_0_RVALID(FringeZynq_io_M_AXI_0_RVALID),
    .io_M_AXI_0_RREADY(FringeZynq_io_M_AXI_0_RREADY),
    .io_M_AXI_0_BID(FringeZynq_io_M_AXI_0_BID),
    .io_M_AXI_0_BVALID(FringeZynq_io_M_AXI_0_BVALID),
    .io_M_AXI_0_BREADY(FringeZynq_io_M_AXI_0_BREADY),
    .io_M_AXI_1_AWID(FringeZynq_io_M_AXI_1_AWID),
    .io_M_AXI_1_AWADDR(FringeZynq_io_M_AXI_1_AWADDR),
    .io_M_AXI_1_AWLEN(FringeZynq_io_M_AXI_1_AWLEN),
    .io_M_AXI_1_AWVALID(FringeZynq_io_M_AXI_1_AWVALID),
    .io_M_AXI_1_AWREADY(FringeZynq_io_M_AXI_1_AWREADY),
    .io_M_AXI_1_ARID(FringeZynq_io_M_AXI_1_ARID),
    .io_M_AXI_1_ARADDR(FringeZynq_io_M_AXI_1_ARADDR),
    .io_M_AXI_1_ARLEN(FringeZynq_io_M_AXI_1_ARLEN),
    .io_M_AXI_1_ARVALID(FringeZynq_io_M_AXI_1_ARVALID),
    .io_M_AXI_1_ARREADY(FringeZynq_io_M_AXI_1_ARREADY),
    .io_M_AXI_1_WDATA(FringeZynq_io_M_AXI_1_WDATA),
    .io_M_AXI_1_WSTRB(FringeZynq_io_M_AXI_1_WSTRB),
    .io_M_AXI_1_WVALID(FringeZynq_io_M_AXI_1_WVALID),
    .io_M_AXI_1_WREADY(FringeZynq_io_M_AXI_1_WREADY),
    .io_M_AXI_1_RID(FringeZynq_io_M_AXI_1_RID),
    .io_M_AXI_1_RDATA(FringeZynq_io_M_AXI_1_RDATA),
    .io_M_AXI_1_RVALID(FringeZynq_io_M_AXI_1_RVALID),
    .io_M_AXI_1_RREADY(FringeZynq_io_M_AXI_1_RREADY),
    .io_M_AXI_1_BID(FringeZynq_io_M_AXI_1_BID),
    .io_M_AXI_1_BVALID(FringeZynq_io_M_AXI_1_BVALID),
    .io_M_AXI_1_BREADY(FringeZynq_io_M_AXI_1_BREADY),
    .io_M_AXI_2_AWID(FringeZynq_io_M_AXI_2_AWID),
    .io_M_AXI_2_AWADDR(FringeZynq_io_M_AXI_2_AWADDR),
    .io_M_AXI_2_AWLEN(FringeZynq_io_M_AXI_2_AWLEN),
    .io_M_AXI_2_AWVALID(FringeZynq_io_M_AXI_2_AWVALID),
    .io_M_AXI_2_AWREADY(FringeZynq_io_M_AXI_2_AWREADY),
    .io_M_AXI_2_ARID(FringeZynq_io_M_AXI_2_ARID),
    .io_M_AXI_2_ARADDR(FringeZynq_io_M_AXI_2_ARADDR),
    .io_M_AXI_2_ARLEN(FringeZynq_io_M_AXI_2_ARLEN),
    .io_M_AXI_2_ARVALID(FringeZynq_io_M_AXI_2_ARVALID),
    .io_M_AXI_2_ARREADY(FringeZynq_io_M_AXI_2_ARREADY),
    .io_M_AXI_2_WDATA(FringeZynq_io_M_AXI_2_WDATA),
    .io_M_AXI_2_WSTRB(FringeZynq_io_M_AXI_2_WSTRB),
    .io_M_AXI_2_WVALID(FringeZynq_io_M_AXI_2_WVALID),
    .io_M_AXI_2_WREADY(FringeZynq_io_M_AXI_2_WREADY),
    .io_M_AXI_2_RID(FringeZynq_io_M_AXI_2_RID),
    .io_M_AXI_2_RDATA(FringeZynq_io_M_AXI_2_RDATA),
    .io_M_AXI_2_RVALID(FringeZynq_io_M_AXI_2_RVALID),
    .io_M_AXI_2_RREADY(FringeZynq_io_M_AXI_2_RREADY),
    .io_M_AXI_2_BID(FringeZynq_io_M_AXI_2_BID),
    .io_M_AXI_2_BVALID(FringeZynq_io_M_AXI_2_BVALID),
    .io_M_AXI_2_BREADY(FringeZynq_io_M_AXI_2_BREADY),
    .io_M_AXI_3_AWID(FringeZynq_io_M_AXI_3_AWID),
    .io_M_AXI_3_AWADDR(FringeZynq_io_M_AXI_3_AWADDR),
    .io_M_AXI_3_AWLEN(FringeZynq_io_M_AXI_3_AWLEN),
    .io_M_AXI_3_AWVALID(FringeZynq_io_M_AXI_3_AWVALID),
    .io_M_AXI_3_AWREADY(FringeZynq_io_M_AXI_3_AWREADY),
    .io_M_AXI_3_ARID(FringeZynq_io_M_AXI_3_ARID),
    .io_M_AXI_3_ARADDR(FringeZynq_io_M_AXI_3_ARADDR),
    .io_M_AXI_3_ARLEN(FringeZynq_io_M_AXI_3_ARLEN),
    .io_M_AXI_3_ARVALID(FringeZynq_io_M_AXI_3_ARVALID),
    .io_M_AXI_3_ARREADY(FringeZynq_io_M_AXI_3_ARREADY),
    .io_M_AXI_3_WDATA(FringeZynq_io_M_AXI_3_WDATA),
    .io_M_AXI_3_WSTRB(FringeZynq_io_M_AXI_3_WSTRB),
    .io_M_AXI_3_WVALID(FringeZynq_io_M_AXI_3_WVALID),
    .io_M_AXI_3_WREADY(FringeZynq_io_M_AXI_3_WREADY),
    .io_M_AXI_3_RID(FringeZynq_io_M_AXI_3_RID),
    .io_M_AXI_3_RDATA(FringeZynq_io_M_AXI_3_RDATA),
    .io_M_AXI_3_RVALID(FringeZynq_io_M_AXI_3_RVALID),
    .io_M_AXI_3_RREADY(FringeZynq_io_M_AXI_3_RREADY),
    .io_M_AXI_3_BID(FringeZynq_io_M_AXI_3_BID),
    .io_M_AXI_3_BVALID(FringeZynq_io_M_AXI_3_BVALID),
    .io_M_AXI_3_BREADY(FringeZynq_io_M_AXI_3_BREADY),
    .io_TOP_AXI_AWADDR(FringeZynq_io_TOP_AXI_AWADDR),
    .io_TOP_AXI_AWLEN(FringeZynq_io_TOP_AXI_AWLEN),
    .io_TOP_AXI_AWVALID(FringeZynq_io_TOP_AXI_AWVALID),
    .io_TOP_AXI_AWREADY(FringeZynq_io_TOP_AXI_AWREADY),
    .io_TOP_AXI_ARID(FringeZynq_io_TOP_AXI_ARID),
    .io_TOP_AXI_ARADDR(FringeZynq_io_TOP_AXI_ARADDR),
    .io_TOP_AXI_ARLEN(FringeZynq_io_TOP_AXI_ARLEN),
    .io_TOP_AXI_ARSIZE(FringeZynq_io_TOP_AXI_ARSIZE),
    .io_TOP_AXI_ARBURST(FringeZynq_io_TOP_AXI_ARBURST),
    .io_TOP_AXI_ARVALID(FringeZynq_io_TOP_AXI_ARVALID),
    .io_TOP_AXI_ARREADY(FringeZynq_io_TOP_AXI_ARREADY),
    .io_TOP_AXI_WDATA(FringeZynq_io_TOP_AXI_WDATA),
    .io_TOP_AXI_WSTRB(FringeZynq_io_TOP_AXI_WSTRB),
    .io_TOP_AXI_WVALID(FringeZynq_io_TOP_AXI_WVALID),
    .io_TOP_AXI_WREADY(FringeZynq_io_TOP_AXI_WREADY),
    .io_TOP_AXI_RVALID(FringeZynq_io_TOP_AXI_RVALID),
    .io_TOP_AXI_RREADY(FringeZynq_io_TOP_AXI_RREADY),
    .io_TOP_AXI_BVALID(FringeZynq_io_TOP_AXI_BVALID),
    .io_TOP_AXI_BREADY(FringeZynq_io_TOP_AXI_BREADY),
    .io_DWIDTH_AXI_AWADDR(FringeZynq_io_DWIDTH_AXI_AWADDR),
    .io_DWIDTH_AXI_AWLEN(FringeZynq_io_DWIDTH_AXI_AWLEN),
    .io_DWIDTH_AXI_AWVALID(FringeZynq_io_DWIDTH_AXI_AWVALID),
    .io_DWIDTH_AXI_AWREADY(FringeZynq_io_DWIDTH_AXI_AWREADY),
    .io_DWIDTH_AXI_ARADDR(FringeZynq_io_DWIDTH_AXI_ARADDR),
    .io_DWIDTH_AXI_ARLEN(FringeZynq_io_DWIDTH_AXI_ARLEN),
    .io_DWIDTH_AXI_ARSIZE(FringeZynq_io_DWIDTH_AXI_ARSIZE),
    .io_DWIDTH_AXI_ARBURST(FringeZynq_io_DWIDTH_AXI_ARBURST),
    .io_DWIDTH_AXI_ARVALID(FringeZynq_io_DWIDTH_AXI_ARVALID),
    .io_DWIDTH_AXI_ARREADY(FringeZynq_io_DWIDTH_AXI_ARREADY),
    .io_DWIDTH_AXI_WDATA(FringeZynq_io_DWIDTH_AXI_WDATA),
    .io_DWIDTH_AXI_WSTRB(FringeZynq_io_DWIDTH_AXI_WSTRB),
    .io_DWIDTH_AXI_WVALID(FringeZynq_io_DWIDTH_AXI_WVALID),
    .io_DWIDTH_AXI_WREADY(FringeZynq_io_DWIDTH_AXI_WREADY),
    .io_DWIDTH_AXI_RVALID(FringeZynq_io_DWIDTH_AXI_RVALID),
    .io_DWIDTH_AXI_RREADY(FringeZynq_io_DWIDTH_AXI_RREADY),
    .io_DWIDTH_AXI_BVALID(FringeZynq_io_DWIDTH_AXI_BVALID),
    .io_DWIDTH_AXI_BREADY(FringeZynq_io_DWIDTH_AXI_BREADY),
    .io_enable(FringeZynq_io_enable),
    .io_done(FringeZynq_io_done),
    .io_reset(FringeZynq_io_reset),
    .io_argIns_0(FringeZynq_io_argIns_0),
    .io_argIns_1(FringeZynq_io_argIns_1),
    .io_argIns_2(FringeZynq_io_argIns_2),
    .io_argOuts_0_valid(FringeZynq_io_argOuts_0_valid),
    .io_argOuts_0_bits(FringeZynq_io_argOuts_0_bits),
    .io_memStreams_loads_3_cmd_ready(FringeZynq_io_memStreams_loads_3_cmd_ready),
    .io_memStreams_loads_3_cmd_valid(FringeZynq_io_memStreams_loads_3_cmd_valid),
    .io_memStreams_loads_3_cmd_bits_addr(FringeZynq_io_memStreams_loads_3_cmd_bits_addr),
    .io_memStreams_loads_3_cmd_bits_isWr(FringeZynq_io_memStreams_loads_3_cmd_bits_isWr),
    .io_memStreams_loads_3_cmd_bits_size(FringeZynq_io_memStreams_loads_3_cmd_bits_size),
    .io_memStreams_loads_3_rdata_ready(FringeZynq_io_memStreams_loads_3_rdata_ready),
    .io_memStreams_loads_3_rdata_valid(FringeZynq_io_memStreams_loads_3_rdata_valid),
    .io_memStreams_loads_3_rdata_bits_0(FringeZynq_io_memStreams_loads_3_rdata_bits_0),
    .io_memStreams_loads_2_cmd_ready(FringeZynq_io_memStreams_loads_2_cmd_ready),
    .io_memStreams_loads_2_cmd_valid(FringeZynq_io_memStreams_loads_2_cmd_valid),
    .io_memStreams_loads_2_cmd_bits_addr(FringeZynq_io_memStreams_loads_2_cmd_bits_addr),
    .io_memStreams_loads_2_cmd_bits_isWr(FringeZynq_io_memStreams_loads_2_cmd_bits_isWr),
    .io_memStreams_loads_2_cmd_bits_size(FringeZynq_io_memStreams_loads_2_cmd_bits_size),
    .io_memStreams_loads_2_rdata_ready(FringeZynq_io_memStreams_loads_2_rdata_ready),
    .io_memStreams_loads_2_rdata_valid(FringeZynq_io_memStreams_loads_2_rdata_valid),
    .io_memStreams_loads_2_rdata_bits_0(FringeZynq_io_memStreams_loads_2_rdata_bits_0),
    .io_memStreams_loads_1_cmd_ready(FringeZynq_io_memStreams_loads_1_cmd_ready),
    .io_memStreams_loads_1_cmd_valid(FringeZynq_io_memStreams_loads_1_cmd_valid),
    .io_memStreams_loads_1_cmd_bits_addr(FringeZynq_io_memStreams_loads_1_cmd_bits_addr),
    .io_memStreams_loads_1_cmd_bits_isWr(FringeZynq_io_memStreams_loads_1_cmd_bits_isWr),
    .io_memStreams_loads_1_cmd_bits_size(FringeZynq_io_memStreams_loads_1_cmd_bits_size),
    .io_memStreams_loads_1_rdata_ready(FringeZynq_io_memStreams_loads_1_rdata_ready),
    .io_memStreams_loads_1_rdata_valid(FringeZynq_io_memStreams_loads_1_rdata_valid),
    .io_memStreams_loads_1_rdata_bits_0(FringeZynq_io_memStreams_loads_1_rdata_bits_0),
    .io_memStreams_loads_0_cmd_ready(FringeZynq_io_memStreams_loads_0_cmd_ready),
    .io_memStreams_loads_0_cmd_valid(FringeZynq_io_memStreams_loads_0_cmd_valid),
    .io_memStreams_loads_0_cmd_bits_addr(FringeZynq_io_memStreams_loads_0_cmd_bits_addr),
    .io_memStreams_loads_0_cmd_bits_isWr(FringeZynq_io_memStreams_loads_0_cmd_bits_isWr),
    .io_memStreams_loads_0_cmd_bits_size(FringeZynq_io_memStreams_loads_0_cmd_bits_size),
    .io_memStreams_loads_0_rdata_ready(FringeZynq_io_memStreams_loads_0_rdata_ready),
    .io_memStreams_loads_0_rdata_valid(FringeZynq_io_memStreams_loads_0_rdata_valid),
    .io_memStreams_loads_0_rdata_bits_0(FringeZynq_io_memStreams_loads_0_rdata_bits_0)
  );
  assign _T_475 = ~ reset;
  assign _T_476 = ~ accel_io_enable;
  assign io_rdata = 1'h0;
  assign io_is_enabled = _T_476;
  assign io_S_AXI_AWREADY = FringeZynq_io_S_AXI_AWREADY;
  assign io_S_AXI_ARREADY = FringeZynq_io_S_AXI_ARREADY;
  assign io_S_AXI_WREADY = FringeZynq_io_S_AXI_WREADY;
  assign io_S_AXI_RDATA = FringeZynq_io_S_AXI_RDATA;
  assign io_S_AXI_RRESP = FringeZynq_io_S_AXI_RRESP;
  assign io_S_AXI_RVALID = FringeZynq_io_S_AXI_RVALID;
  assign io_S_AXI_BRESP = FringeZynq_io_S_AXI_BRESP;
  assign io_S_AXI_BVALID = FringeZynq_io_S_AXI_BVALID;
  assign io_M_AXI_0_AWID = FringeZynq_io_M_AXI_0_AWID;
  assign io_M_AXI_0_AWUSER = 32'h0;
  assign io_M_AXI_0_AWADDR = FringeZynq_io_M_AXI_0_AWADDR;
  assign io_M_AXI_0_AWLEN = FringeZynq_io_M_AXI_0_AWLEN;
  assign io_M_AXI_0_AWSIZE = 3'h6;
  assign io_M_AXI_0_AWBURST = 2'h1;
  assign io_M_AXI_0_AWLOCK = 1'h0;
  assign io_M_AXI_0_AWCACHE = 4'h3;
  assign io_M_AXI_0_AWPROT = 3'h0;
  assign io_M_AXI_0_AWQOS = 4'h0;
  assign io_M_AXI_0_AWVALID = FringeZynq_io_M_AXI_0_AWVALID;
  assign io_M_AXI_0_ARID = FringeZynq_io_M_AXI_0_ARID;
  assign io_M_AXI_0_ARUSER = 32'h0;
  assign io_M_AXI_0_ARADDR = FringeZynq_io_M_AXI_0_ARADDR;
  assign io_M_AXI_0_ARLEN = FringeZynq_io_M_AXI_0_ARLEN;
  assign io_M_AXI_0_ARSIZE = 3'h6;
  assign io_M_AXI_0_ARBURST = 2'h1;
  assign io_M_AXI_0_ARLOCK = 1'h0;
  assign io_M_AXI_0_ARCACHE = 4'h3;
  assign io_M_AXI_0_ARPROT = 3'h0;
  assign io_M_AXI_0_ARQOS = 4'h0;
  assign io_M_AXI_0_ARVALID = FringeZynq_io_M_AXI_0_ARVALID;
  assign io_M_AXI_0_WDATA = FringeZynq_io_M_AXI_0_WDATA;
  assign io_M_AXI_0_WSTRB = FringeZynq_io_M_AXI_0_WSTRB;
  assign io_M_AXI_0_WLAST = 1'h0;
  assign io_M_AXI_0_WVALID = FringeZynq_io_M_AXI_0_WVALID;
  assign io_M_AXI_0_RREADY = FringeZynq_io_M_AXI_0_RREADY;
  assign io_M_AXI_0_BREADY = FringeZynq_io_M_AXI_0_BREADY;
  assign io_M_AXI_1_AWID = FringeZynq_io_M_AXI_1_AWID;
  assign io_M_AXI_1_AWUSER = 32'h0;
  assign io_M_AXI_1_AWADDR = FringeZynq_io_M_AXI_1_AWADDR;
  assign io_M_AXI_1_AWLEN = FringeZynq_io_M_AXI_1_AWLEN;
  assign io_M_AXI_1_AWSIZE = 3'h6;
  assign io_M_AXI_1_AWBURST = 2'h1;
  assign io_M_AXI_1_AWLOCK = 1'h0;
  assign io_M_AXI_1_AWCACHE = 4'h3;
  assign io_M_AXI_1_AWPROT = 3'h0;
  assign io_M_AXI_1_AWQOS = 4'h0;
  assign io_M_AXI_1_AWVALID = FringeZynq_io_M_AXI_1_AWVALID;
  assign io_M_AXI_1_ARID = FringeZynq_io_M_AXI_1_ARID;
  assign io_M_AXI_1_ARUSER = 32'h0;
  assign io_M_AXI_1_ARADDR = FringeZynq_io_M_AXI_1_ARADDR;
  assign io_M_AXI_1_ARLEN = FringeZynq_io_M_AXI_1_ARLEN;
  assign io_M_AXI_1_ARSIZE = 3'h6;
  assign io_M_AXI_1_ARBURST = 2'h1;
  assign io_M_AXI_1_ARLOCK = 1'h0;
  assign io_M_AXI_1_ARCACHE = 4'h3;
  assign io_M_AXI_1_ARPROT = 3'h0;
  assign io_M_AXI_1_ARQOS = 4'h0;
  assign io_M_AXI_1_ARVALID = FringeZynq_io_M_AXI_1_ARVALID;
  assign io_M_AXI_1_WDATA = FringeZynq_io_M_AXI_1_WDATA;
  assign io_M_AXI_1_WSTRB = FringeZynq_io_M_AXI_1_WSTRB;
  assign io_M_AXI_1_WLAST = 1'h0;
  assign io_M_AXI_1_WVALID = FringeZynq_io_M_AXI_1_WVALID;
  assign io_M_AXI_1_RREADY = FringeZynq_io_M_AXI_1_RREADY;
  assign io_M_AXI_1_BREADY = FringeZynq_io_M_AXI_1_BREADY;
  assign io_M_AXI_2_AWID = FringeZynq_io_M_AXI_2_AWID;
  assign io_M_AXI_2_AWUSER = 32'h0;
  assign io_M_AXI_2_AWADDR = FringeZynq_io_M_AXI_2_AWADDR;
  assign io_M_AXI_2_AWLEN = FringeZynq_io_M_AXI_2_AWLEN;
  assign io_M_AXI_2_AWSIZE = 3'h6;
  assign io_M_AXI_2_AWBURST = 2'h1;
  assign io_M_AXI_2_AWLOCK = 1'h0;
  assign io_M_AXI_2_AWCACHE = 4'h3;
  assign io_M_AXI_2_AWPROT = 3'h0;
  assign io_M_AXI_2_AWQOS = 4'h0;
  assign io_M_AXI_2_AWVALID = FringeZynq_io_M_AXI_2_AWVALID;
  assign io_M_AXI_2_ARID = FringeZynq_io_M_AXI_2_ARID;
  assign io_M_AXI_2_ARUSER = 32'h0;
  assign io_M_AXI_2_ARADDR = FringeZynq_io_M_AXI_2_ARADDR;
  assign io_M_AXI_2_ARLEN = FringeZynq_io_M_AXI_2_ARLEN;
  assign io_M_AXI_2_ARSIZE = 3'h6;
  assign io_M_AXI_2_ARBURST = 2'h1;
  assign io_M_AXI_2_ARLOCK = 1'h0;
  assign io_M_AXI_2_ARCACHE = 4'h3;
  assign io_M_AXI_2_ARPROT = 3'h0;
  assign io_M_AXI_2_ARQOS = 4'h0;
  assign io_M_AXI_2_ARVALID = FringeZynq_io_M_AXI_2_ARVALID;
  assign io_M_AXI_2_WDATA = FringeZynq_io_M_AXI_2_WDATA;
  assign io_M_AXI_2_WSTRB = FringeZynq_io_M_AXI_2_WSTRB;
  assign io_M_AXI_2_WLAST = 1'h0;
  assign io_M_AXI_2_WVALID = FringeZynq_io_M_AXI_2_WVALID;
  assign io_M_AXI_2_RREADY = FringeZynq_io_M_AXI_2_RREADY;
  assign io_M_AXI_2_BREADY = FringeZynq_io_M_AXI_2_BREADY;
  assign io_M_AXI_3_AWID = FringeZynq_io_M_AXI_3_AWID;
  assign io_M_AXI_3_AWUSER = 32'h0;
  assign io_M_AXI_3_AWADDR = FringeZynq_io_M_AXI_3_AWADDR;
  assign io_M_AXI_3_AWLEN = FringeZynq_io_M_AXI_3_AWLEN;
  assign io_M_AXI_3_AWSIZE = 3'h6;
  assign io_M_AXI_3_AWBURST = 2'h1;
  assign io_M_AXI_3_AWLOCK = 1'h0;
  assign io_M_AXI_3_AWCACHE = 4'h3;
  assign io_M_AXI_3_AWPROT = 3'h0;
  assign io_M_AXI_3_AWQOS = 4'h0;
  assign io_M_AXI_3_AWVALID = FringeZynq_io_M_AXI_3_AWVALID;
  assign io_M_AXI_3_ARID = FringeZynq_io_M_AXI_3_ARID;
  assign io_M_AXI_3_ARUSER = 32'h0;
  assign io_M_AXI_3_ARADDR = FringeZynq_io_M_AXI_3_ARADDR;
  assign io_M_AXI_3_ARLEN = FringeZynq_io_M_AXI_3_ARLEN;
  assign io_M_AXI_3_ARSIZE = 3'h6;
  assign io_M_AXI_3_ARBURST = 2'h1;
  assign io_M_AXI_3_ARLOCK = 1'h0;
  assign io_M_AXI_3_ARCACHE = 4'h3;
  assign io_M_AXI_3_ARPROT = 3'h0;
  assign io_M_AXI_3_ARQOS = 4'h0;
  assign io_M_AXI_3_ARVALID = FringeZynq_io_M_AXI_3_ARVALID;
  assign io_M_AXI_3_WDATA = FringeZynq_io_M_AXI_3_WDATA;
  assign io_M_AXI_3_WSTRB = FringeZynq_io_M_AXI_3_WSTRB;
  assign io_M_AXI_3_WLAST = 1'h0;
  assign io_M_AXI_3_WVALID = FringeZynq_io_M_AXI_3_WVALID;
  assign io_M_AXI_3_RREADY = FringeZynq_io_M_AXI_3_RREADY;
  assign io_M_AXI_3_BREADY = FringeZynq_io_M_AXI_3_BREADY;
  assign accel_io_enable = FringeZynq_io_enable;
  assign accel_io_memStreams_loads_3_cmd_ready = FringeZynq_io_memStreams_loads_3_cmd_ready;
  assign accel_io_memStreams_loads_3_rdata_valid = FringeZynq_io_memStreams_loads_3_rdata_valid;
  assign accel_io_memStreams_loads_3_rdata_bits_0 = FringeZynq_io_memStreams_loads_3_rdata_bits_0;
  assign accel_io_memStreams_loads_2_cmd_ready = FringeZynq_io_memStreams_loads_2_cmd_ready;
  assign accel_io_memStreams_loads_2_rdata_valid = FringeZynq_io_memStreams_loads_2_rdata_valid;
  assign accel_io_memStreams_loads_2_rdata_bits_0 = FringeZynq_io_memStreams_loads_2_rdata_bits_0;
  assign accel_io_memStreams_loads_1_cmd_ready = FringeZynq_io_memStreams_loads_1_cmd_ready;
  assign accel_io_memStreams_loads_1_rdata_valid = FringeZynq_io_memStreams_loads_1_rdata_valid;
  assign accel_io_memStreams_loads_1_rdata_bits_0 = FringeZynq_io_memStreams_loads_1_rdata_bits_0;
  assign accel_io_memStreams_loads_0_cmd_ready = FringeZynq_io_memStreams_loads_0_cmd_ready;
  assign accel_io_memStreams_loads_0_rdata_valid = FringeZynq_io_memStreams_loads_0_rdata_valid;
  assign accel_io_memStreams_loads_0_rdata_bits_0 = FringeZynq_io_memStreams_loads_0_rdata_bits_0;
  assign accel_io_argIns_0 = FringeZynq_io_argIns_0;
  assign accel_io_argIns_1 = FringeZynq_io_argIns_1;
  assign accel_io_argIns_2 = FringeZynq_io_argIns_2;
  assign accel_clock = clock;
  assign accel_reset = FringeZynq_io_reset;
  assign FringeZynq_io_S_AXI_AWADDR = io_S_AXI_AWADDR;
  assign FringeZynq_io_S_AXI_AWPROT = io_S_AXI_AWPROT;
  assign FringeZynq_io_S_AXI_AWVALID = io_S_AXI_AWVALID;
  assign FringeZynq_io_S_AXI_ARADDR = io_S_AXI_ARADDR;
  assign FringeZynq_io_S_AXI_ARPROT = io_S_AXI_ARPROT;
  assign FringeZynq_io_S_AXI_ARVALID = io_S_AXI_ARVALID;
  assign FringeZynq_io_S_AXI_WDATA = io_S_AXI_WDATA;
  assign FringeZynq_io_S_AXI_WSTRB = io_S_AXI_WSTRB;
  assign FringeZynq_io_S_AXI_WVALID = io_S_AXI_WVALID;
  assign FringeZynq_io_S_AXI_RREADY = io_S_AXI_RREADY;
  assign FringeZynq_io_S_AXI_BREADY = io_S_AXI_BREADY;
  assign FringeZynq_io_M_AXI_0_AWREADY = io_M_AXI_0_AWREADY;
  assign FringeZynq_io_M_AXI_0_ARREADY = io_M_AXI_0_ARREADY;
  assign FringeZynq_io_M_AXI_0_WREADY = io_M_AXI_0_WREADY;
  assign FringeZynq_io_M_AXI_0_RID = io_M_AXI_0_RID;
  assign FringeZynq_io_M_AXI_0_RDATA = io_M_AXI_0_RDATA;
  assign FringeZynq_io_M_AXI_0_RVALID = io_M_AXI_0_RVALID;
  assign FringeZynq_io_M_AXI_0_BID = io_M_AXI_0_BID;
  assign FringeZynq_io_M_AXI_0_BVALID = io_M_AXI_0_BVALID;
  assign FringeZynq_io_M_AXI_1_AWREADY = io_M_AXI_1_AWREADY;
  assign FringeZynq_io_M_AXI_1_ARREADY = io_M_AXI_1_ARREADY;
  assign FringeZynq_io_M_AXI_1_WREADY = io_M_AXI_1_WREADY;
  assign FringeZynq_io_M_AXI_1_RID = io_M_AXI_1_RID;
  assign FringeZynq_io_M_AXI_1_RDATA = io_M_AXI_1_RDATA;
  assign FringeZynq_io_M_AXI_1_RVALID = io_M_AXI_1_RVALID;
  assign FringeZynq_io_M_AXI_1_BID = io_M_AXI_1_BID;
  assign FringeZynq_io_M_AXI_1_BVALID = io_M_AXI_1_BVALID;
  assign FringeZynq_io_M_AXI_2_AWREADY = io_M_AXI_2_AWREADY;
  assign FringeZynq_io_M_AXI_2_ARREADY = io_M_AXI_2_ARREADY;
  assign FringeZynq_io_M_AXI_2_WREADY = io_M_AXI_2_WREADY;
  assign FringeZynq_io_M_AXI_2_RID = io_M_AXI_2_RID;
  assign FringeZynq_io_M_AXI_2_RDATA = io_M_AXI_2_RDATA;
  assign FringeZynq_io_M_AXI_2_RVALID = io_M_AXI_2_RVALID;
  assign FringeZynq_io_M_AXI_2_BID = io_M_AXI_2_BID;
  assign FringeZynq_io_M_AXI_2_BVALID = io_M_AXI_2_BVALID;
  assign FringeZynq_io_M_AXI_3_AWREADY = io_M_AXI_3_AWREADY;
  assign FringeZynq_io_M_AXI_3_ARREADY = io_M_AXI_3_ARREADY;
  assign FringeZynq_io_M_AXI_3_WREADY = io_M_AXI_3_WREADY;
  assign FringeZynq_io_M_AXI_3_RID = io_M_AXI_3_RID;
  assign FringeZynq_io_M_AXI_3_RDATA = io_M_AXI_3_RDATA;
  assign FringeZynq_io_M_AXI_3_RVALID = io_M_AXI_3_RVALID;
  assign FringeZynq_io_M_AXI_3_BID = io_M_AXI_3_BID;
  assign FringeZynq_io_M_AXI_3_BVALID = io_M_AXI_3_BVALID;
  assign FringeZynq_io_TOP_AXI_AWADDR = io_TOP_AXI_AWADDR;
  assign FringeZynq_io_TOP_AXI_AWLEN = io_TOP_AXI_AWLEN;
  assign FringeZynq_io_TOP_AXI_AWVALID = io_TOP_AXI_AWVALID;
  assign FringeZynq_io_TOP_AXI_AWREADY = io_TOP_AXI_AWREADY;
  assign FringeZynq_io_TOP_AXI_ARID = io_TOP_AXI_ARID;
  assign FringeZynq_io_TOP_AXI_ARADDR = io_TOP_AXI_ARADDR;
  assign FringeZynq_io_TOP_AXI_ARLEN = io_TOP_AXI_ARLEN;
  assign FringeZynq_io_TOP_AXI_ARSIZE = io_TOP_AXI_ARSIZE;
  assign FringeZynq_io_TOP_AXI_ARBURST = io_TOP_AXI_ARBURST;
  assign FringeZynq_io_TOP_AXI_ARVALID = io_TOP_AXI_ARVALID;
  assign FringeZynq_io_TOP_AXI_ARREADY = io_TOP_AXI_ARREADY;
  assign FringeZynq_io_TOP_AXI_WDATA = io_TOP_AXI_WDATA;
  assign FringeZynq_io_TOP_AXI_WSTRB = io_TOP_AXI_WSTRB;
  assign FringeZynq_io_TOP_AXI_WVALID = io_TOP_AXI_WVALID;
  assign FringeZynq_io_TOP_AXI_WREADY = io_TOP_AXI_WREADY;
  assign FringeZynq_io_TOP_AXI_RVALID = io_TOP_AXI_RVALID;
  assign FringeZynq_io_TOP_AXI_RREADY = io_TOP_AXI_RREADY;
  assign FringeZynq_io_TOP_AXI_BVALID = io_TOP_AXI_BVALID;
  assign FringeZynq_io_TOP_AXI_BREADY = io_TOP_AXI_BREADY;
  assign FringeZynq_io_DWIDTH_AXI_AWADDR = io_DWIDTH_AXI_AWADDR;
  assign FringeZynq_io_DWIDTH_AXI_AWLEN = io_DWIDTH_AXI_AWLEN;
  assign FringeZynq_io_DWIDTH_AXI_AWVALID = io_DWIDTH_AXI_AWVALID;
  assign FringeZynq_io_DWIDTH_AXI_AWREADY = io_DWIDTH_AXI_AWREADY;
  assign FringeZynq_io_DWIDTH_AXI_ARADDR = io_DWIDTH_AXI_ARADDR;
  assign FringeZynq_io_DWIDTH_AXI_ARLEN = io_DWIDTH_AXI_ARLEN;
  assign FringeZynq_io_DWIDTH_AXI_ARSIZE = io_DWIDTH_AXI_ARSIZE;
  assign FringeZynq_io_DWIDTH_AXI_ARBURST = io_DWIDTH_AXI_ARBURST;
  assign FringeZynq_io_DWIDTH_AXI_ARVALID = io_DWIDTH_AXI_ARVALID;
  assign FringeZynq_io_DWIDTH_AXI_ARREADY = io_DWIDTH_AXI_ARREADY;
  assign FringeZynq_io_DWIDTH_AXI_WDATA = io_DWIDTH_AXI_WDATA;
  assign FringeZynq_io_DWIDTH_AXI_WSTRB = io_DWIDTH_AXI_WSTRB;
  assign FringeZynq_io_DWIDTH_AXI_WVALID = io_DWIDTH_AXI_WVALID;
  assign FringeZynq_io_DWIDTH_AXI_WREADY = io_DWIDTH_AXI_WREADY;
  assign FringeZynq_io_DWIDTH_AXI_RVALID = io_DWIDTH_AXI_RVALID;
  assign FringeZynq_io_DWIDTH_AXI_RREADY = io_DWIDTH_AXI_RREADY;
  assign FringeZynq_io_DWIDTH_AXI_BVALID = io_DWIDTH_AXI_BVALID;
  assign FringeZynq_io_DWIDTH_AXI_BREADY = io_DWIDTH_AXI_BREADY;
  assign FringeZynq_io_done = accel_io_done;
  assign FringeZynq_io_argOuts_0_valid = accel_io_argOuts_0_valid;
  assign FringeZynq_io_argOuts_0_bits = accel_io_argOuts_0_bits;
  assign FringeZynq_io_memStreams_loads_3_cmd_valid = accel_io_memStreams_loads_3_cmd_valid;
  assign FringeZynq_io_memStreams_loads_3_cmd_bits_addr = accel_io_memStreams_loads_3_cmd_bits_addr;
  assign FringeZynq_io_memStreams_loads_3_cmd_bits_isWr = accel_io_memStreams_loads_3_cmd_bits_isWr;
  assign FringeZynq_io_memStreams_loads_3_cmd_bits_size = accel_io_memStreams_loads_3_cmd_bits_size;
  assign FringeZynq_io_memStreams_loads_3_rdata_ready = accel_io_memStreams_loads_3_rdata_ready;
  assign FringeZynq_io_memStreams_loads_2_cmd_valid = accel_io_memStreams_loads_2_cmd_valid;
  assign FringeZynq_io_memStreams_loads_2_cmd_bits_addr = accel_io_memStreams_loads_2_cmd_bits_addr;
  assign FringeZynq_io_memStreams_loads_2_cmd_bits_isWr = accel_io_memStreams_loads_2_cmd_bits_isWr;
  assign FringeZynq_io_memStreams_loads_2_cmd_bits_size = accel_io_memStreams_loads_2_cmd_bits_size;
  assign FringeZynq_io_memStreams_loads_2_rdata_ready = accel_io_memStreams_loads_2_rdata_ready;
  assign FringeZynq_io_memStreams_loads_1_cmd_valid = accel_io_memStreams_loads_1_cmd_valid;
  assign FringeZynq_io_memStreams_loads_1_cmd_bits_addr = accel_io_memStreams_loads_1_cmd_bits_addr;
  assign FringeZynq_io_memStreams_loads_1_cmd_bits_isWr = accel_io_memStreams_loads_1_cmd_bits_isWr;
  assign FringeZynq_io_memStreams_loads_1_cmd_bits_size = accel_io_memStreams_loads_1_cmd_bits_size;
  assign FringeZynq_io_memStreams_loads_1_rdata_ready = accel_io_memStreams_loads_1_rdata_ready;
  assign FringeZynq_io_memStreams_loads_0_cmd_valid = accel_io_memStreams_loads_0_cmd_valid;
  assign FringeZynq_io_memStreams_loads_0_cmd_bits_addr = accel_io_memStreams_loads_0_cmd_bits_addr;
  assign FringeZynq_io_memStreams_loads_0_cmd_bits_isWr = accel_io_memStreams_loads_0_cmd_bits_isWr;
  assign FringeZynq_io_memStreams_loads_0_cmd_bits_size = accel_io_memStreams_loads_0_cmd_bits_size;
  assign FringeZynq_io_memStreams_loads_0_rdata_ready = accel_io_memStreams_loads_0_rdata_ready;
  assign FringeZynq_clock = clock;
  assign FringeZynq_reset = _T_475;
endmodule
module SRAMVerilogAWS
#(
    parameter WORDS = 1024,
    parameter AWIDTH = 10,
    parameter DWIDTH = 32)
(
    input clk,
    input [AWIDTH-1:0] raddr,
    input [AWIDTH-1:0] waddr,
    input raddrEn,
    input waddrEn,
    input wen,
    input [DWIDTH-1:0] wdata,
    input flow,
    output reg [DWIDTH-1:0] rdata
);

    reg [DWIDTH-1:0] mem [0:WORDS-1];

    always @(posedge clk) begin
      if (wen) mem[waddr] <= wdata;
      if (flow) rdata <= mem[raddr];
    end

endmodule
